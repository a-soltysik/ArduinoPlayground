PK   <?X���A  F4    cirkitFile.json�[o#Wv��J�ygׅ�~g&�&c����� Jdq�Y�P�/1����b_(�(���5�C8c��ŏ��v�*���Ѯ���],��v�S���loG����ov����G�����v��.��k>�������Ў�wm����mEY��d^��M}=��Y;�_7��IeU1���4i��o��ͻ��+XX!k��
iQ��
iQ��
iQ��
iQ��
i1	3D�bf�*��,�UH�y�!��5�2,�E�R��/�a�,/�a�,/�a�,/�a�,/�a�,/�a�,/�a�,���r���m{�_�괴yZ�'ӪWi�_Ϛzܔ6+��ӶY�(�	�u���ݰD��>�@`�� Nq�s�x�.�e;,�)�e;,�)�e;,�)�e;,�)��RUF��x�/�%?,�U�c?lnw�]���\`�a{��6�_Ƿ�?F��t$~)㇐�D�����%2E�������1����"~Kd��1 ,�)��a�L��a�L���H�*^;��"^;��"^;��"^;���N��U�v�%2E�v�%2E�v�%2E�v�%2E�v�%Ң��ΰD���ΰD���ΰD���ΰD���ΰD� ~e���:^;��"^;��"^;��"^;�i1��ΰD���ΰD���Ξ���B��U��;R�/2.��tA1��Y��Ō2�w#錥3�.-
ֻ���3�.-Jֻ���3�.�ֻ���3�.���լw(��t�L��n�z��K�Sֻ)�Jg,]Z�X�f�w(��ti1g���ޡt���M���1z�n0��|~;)��.�x����	��3��o���S�g0��|�'��`>�m�N,��|~�7��8X>���Vu�?8u�|��M��p�`�����p�`����	�f8�|�����p�`�����/�Op�(��Q����3��g�������3����������3��g.������3���\������3��g|������3���T3Ŀ��}侫�9�/��/���'�/%_X>��|J�_X>��|2"�_X>��|%�}�}�_J8��p|a��󩫰p|a���I��p|a����°p|a���ΰp|a���)ڰ��',��|>�������g0�O������g0�O�����g0��"�����g0�7Q���'��3E��Q������g0�7������g0��܀����g0�7�����g0��9�����g0�7ha��������e`�������Mq`��������|`������獈`�������-�`�����lu8�p��������m�`��������`��������`�������M�X�&p�`����l�p�`����r�p�`����m�N��Z�������O���������Oۆ�������Ou�������O[c6�aw�uۆny��҆n{��Ɇ7����rr��G�ٵŦV6�v9���?I�mm�xڔ�tU���4[X������շŦ�<����������ޒUC����n�qzK=xGo����'3���rl����O��O9/WMS5�T,��3��6����E��?�L�:͗u9Nv�d���xV�i<k�d�i[5�z�_����~���?�E��������i����}����f��/|>�S���,qf�P�c0D�P��1D�P��2D�P�`:C	u˧3D�P��:C	uK�3D�P��:C	uˮ3D�P��/T"��͕m�nV�)��%�	�݆oJ)uW( &�~V�)��]I���nX���KYiަ4k�LX/�:N)�x��f�?S���o���V�)��j�V���SJ���!&����k)M�A&��X���C�	��%V�)��:�V�K��SJ�5�!&���X���CLX/�:N)�n���:^bu�R:��1au���8�tX�b��x��qJ�<��]�.�cu���8�tX9b��x��qJ鰪<Ą��
���a�y����X����CLX��:N)V����_7��7�:^cu�R:�i1au���8�tX�b�����R�����:>���9���ݜ\����ؕ��"��+���\\c5	�IXSoz\�U�j��[�W}U���5�V��UA_�&aM���qU�W�IXSo�{\�U�jִ8�-����*XM�=pU�W�IX���
��`5	���	�cZ�����oE�K�4��4��4�KBkZ��\�&}IhMC���k��$0	�ih�����&�5��a�x�IbZ���\���4&�5��)�x�IdZ�������T&�5��������eZ���\%���\&�5�Ϲ�x+�EL���&��\Vhr���4�>N�&�IhMC�s�4�jr���4�>'Q�&�IhMC�s+5�jr���4�>GT�&�IhMC�s]5���q����%L(5����2	�ih}��[M.�К���Pk���2	�ih}.��[�݊��5����R��$������o5�LBkZ�1��V��$����^	o5�LBkZ����V��$�����o5��IhMC�=8$�V�\&�5���x��eZ��zO���\&�5��v�x��eZ��z�����d��d�\VirY��eZ��z� ���\&�5��>�x��eZ��z'���\&�5����x��eZ��zO-���&�IhMC��4�jr���4���L�&�IhMC��4�jr���4��sN�&�IhMC��4ފ�|��|hrY��e�&�IhMC�5�jr���4�ޓQ�&�IhMC�%5�jr���4��#S��D��$����^�o5�LBkZ�Y��V��$�v��%��t���4�r���Ѕ��3�����=P�Lw�*g�QT9�Az�ʙ��CG4x��{n�ס2��=���Pf�[�t�L7���O��0����uJe�z�(>�~�P�n�>*sŽ�	��0���Z�Ce�Q|n�š2�(>���У.3�ϭ�Uf>��Ԯ�c[�f~�T�s�r:^���j�X���g5�0,�.Ry��0��4_��8�u����Yݦ�)���m���y_.Ry֗�T���"�g}�Z٬��t��R>�.�ag�xڔ�tU���4{ޗ�T��x�Y췋�}�oG��*;|��m�����o����a�@� ��~�AB�}!��R�j"H(u		!��R��"H(u�!��R�"H(u�!���!�2%���\���a��RJ��0a�۰�M)����	�߆pJ).\0LX7��SJ�pI�a��x��qJ).�0L��7w�����R:\�b��:^`u�RJ��mV���SJ�p�a��x��qJ)�P2q��%V�)%��1qWR�K)X/�:N)y�	��%V�)%���1au���8��=&0&��WX����Ƅ��
�㔒ϡǘ�k��Eq��WX��|�3Ƅ��
�㔒ϭŘ�:^au�R��O?X��:N)��A�	��5V�)%���1q�nr?obu���8��s�0&���X��|Ƅ��	V�)%�3�1au|���sJ��?���Ъ�i
��IXM��
_{Sk�&aM�޼Z�U�jִ��:�UA_�&a͹K�k�� �$��<H�k�� �$��E�k�� �$�i��m@���*XM���*諂�$�i��i@���*XM���k��&qIhMC��6k��.Q���.�/�$/	�ih�^s����%�5��3��V��$����{�5�jR���4�>�A�&�IhMC�s14�jҘ��4�>�D�&�IhMC�sc4�jR���4�>�G�Â&�IhMC�s�4�jr���4�>�J��1�Ob�\VhrY��eZ���8���\&�5����x��eZ����D���\&�5�ϭ�x��eZ���Q���\&�5��u�x��eZ����]͍I�\&�5��=�x��eZ���j���\&�5���x+�[Qt��&���\Vjr���4�>7_�&�IhMC�=4�jr���4��+A�&�IhMC�=4�jr���4�޻B�&�IhMC�=8$�V�\&�5���x��eZ��zO���\&�5��v�x��eZ��z�����d��d�\VirY��eZ��z� ���\&�5��>�x��eZ��z'���\&�5����x��eZ��zO-���&�IhMC��4�jr���4���L�&�IhMC��4�jr���4��sN�&�IhMC��4ފ�|��|hrY��e�&�IhMC�5�jr���4�ޓQ�&�IhMC�%5�jr���4��#S��D��$����^�o5�LBkZ�Y��V��$�v��u��t��r�7����3}����=P�L��*g�[T9ӏz�ʙ�U��|:��ˌ�s���a�﹥U��0#���Ce�1|n�С2�(>��P�3���*�Ce�Q|n-ȡ2�(>���Pf�[�p�Q���V�*3��lj�˱�V3?W*�R9/WMS5�T,������T�gw��T�ݟ&U��˺'�n���z<��4�5E����[=��E*��r�ʳ�\��/S+�u����U���E7�O������u�f��r�ʱ/����_,�7��b��e�zr5�y�k�n�e�Zln�ݪݍ^�y9$��I~w�&�v:���Ek�>�y�B��?��~{�"��6���$��)��W�9��5��*F�ʃ�^7�l�c����n~�הc	���r�C������>v�۟��]=v�x�!����9���p�z���9zſP� P �2�8�!C>�uL(�O;v�)����42x*����<Z=�rn����@��T��/�_sZt�θ�{��=7P~w�g\���~b�����v���7�v������� ��o�����o���Q�C��%��a��e� EX�p�0H�Hݏ�A��D�~�R�%R�cn�",����a�����K���� EX"~̎�-�z���иF:�� j�E4��wD9�:j@!�k��=	Q��PL��pWDz�O��$��c@y�k��m'�X�8[%NW�j[ �6��7�D9�j[ �6����D9�j��;s���.�A2�߸F:��W���@�k���EQ�ږ@��kx�Y���%Pm���� �m	T۸���8��Z�5��-��V@=�kx+?���PO��"� ��\�zZ�4��m� ��V@=�kx�'���PO��V�i ��5PO�ޮ� �i�Ӹ��A8�_�����zZ�4��( ���@=�kx�������5|�<���	PO���k��9��|��KO)"o0��q���A����3�/-z]8=�?��`���u����X>���u���k?��,��|�t���b.�yY>���i�_��\��|�E�c�����̗��p���g0_Z�:�qz�,��|~�#}͞�Mh4�߮I{��<��9�t�*�xHG��o��=��Lh4a*�xHG��oO�=�S	Lh4��ZM{H'��hB�-���N'0�ф~K;�!�P`B�	�v|�C:���F���B5�S`B�	}��!�S`B�	}��!��	��	�S
:�tN�	�&��1��tN�	�&�=��tN�	�&�II��tN�	�&�	U��tN�	�&��_��tN�	�&|؂�����������Aǖ��-0�ф>c����-0�ф>ۑ���-0�ф>S�����ۋ�-%[J:���F�Y�C:���F��^�C:���F��d�C:���F��j�C:���F��p�C����hB��{X�9&4��g���9&4�л��9&4��; ��9&4�л7��S�)tN��R�9&4�лf��9&4��;~��9&4�л���9&4��;���9&4�л���tN�	�&�7��tN�	�&��<��tN�	�&��B��tN�	�&��H��tN�	�&�N���$z|=�Sj:��tN�	�&�NZ��tN�	�&�.`��tN�	�&�f��tN�	�&��k��:���Fz�8�C:���Fz�;�C:�������{�.�ܾ�qp���Ϋ��uL�}�����{Jn��,:p�^GЁ��:y?���܆
D�`ɴ��Q�_�l��#k�D���6|Y�P�S�q�_Ak���O/z6T�����(�!5|=��@����W*���%��
<1N瓙M�z9��j�g(e>C)���i�f���<=uFq������_���|R�i���q��&X�ǳ�M�YS$[O۪��S������m���h�'>�E��?��/\������j�Uf��ĳ���%~ɨ�~3�Ñ����uӏu�w����g�__�ݺ�+�_j�Z�������7ߠ[Ͻ�-�N۷(|�·(|�·(|�·(|�ҷ�{ڻ����>~��/��/��n�.[p��ݻ��d���_?� �����v��t���E�ޅ O'�]�`�OXD�/B��vK&���Qh�Eo!�Qu��º:=ڏ��/��Ms�����ߏF�������� �Sŧ���S姧��Sէ������,�|�ܮ������=���I�(���o�j~�Ϭ�-��M���W�/x�/_��_����ߺ���m?�����?~����o3�p��mn}��m~���٫�O�ͽ��g7k�u��v�iG����o���g���uss��'�������M��]�?��]�+�>cg�ln���r�kwO��d����n���a{��o�ه7�"����լ�����N�m~i�ZV�u����xZ��I��x��Qu=��U�c��?���NҮF� �on����W��n�U�����kov˛��W�I��Uu��O�����?���36/^�_��N���?S?S?cG�̎�{z���������X����G��{_}y���~��ϔ'�ؗg��6ɾ��͎�i����3��3���H��?fGOL�����/��>?���������_m�_���^��R.Tѝ٬;i����U���o������޷ɟ߫���Y5/�ʫjR���?I��R��˲^'/�y����*'�|6j��dy����uy��~�i�%�{�>8�]�?�������y9�tX�2H��aV}v�D��G$�HrC�x5�:�_�Ru4 ?}��xQZ�h<��"�����ȼ�\�N_�yl}���u^M��X<����zr������w���0\�����������|��Ng�y�N��z>}��\�?8=�Wu�L��q��g5�IZ�Ӫ�q9�'FUդ�q���(�_tzTwG�t8��'�prU�>�����g����U7J����,�W��r5�N�_�rq���ϛ����R}�}���{�d��<��閿>P��=��}���K\�n������i�����yf��mv�f�{;z�v�'����M�vt�6��f��ns��{��%:��v��V�*E'�k~�e͂��~�nn��5����oo߾y~���;��n���G_���ߝ�~������E�գ/�<���s��t��wߎ>�!7x���:�N.#=7��������o��������'��G��퉯�ţI����C��^T?�xy�W���'����ǿ�|hN�)��?u�|QV�mO�ۿ_;�..ءO^5���<zUe/yY���p��)�Zx��S���W�u�Ş=�v�p)//��wz��ΝOt����q��)��Z/���S���El�(��7���~8��$��_h1}8�.{٤~|�u�]����(�h������o;�mr���)������������|����}���wG�PK   <?X�����  �  /   images/37b7845a-1f46-4418-9ae8-cf8221840334.png�5�PNG

   IHDR   d   s   n1�w   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  WIDATx��k�E�k�Ǡ�y��vD��.��"�btW�&�,����1�F��Ȣ�5*j| �� ��ET��(�DQy�֯�3).]}������?��̝��U��s�S��*O����?�r�.�ui��6]��r�.k�SO=U%��z���_��֥�.�tY��m�̑�|��!���]*��Z��GUC�]>T飳�$=����O�ٺ�E�)|�d�u�)�x��B�Q�;]��ɰ�A��T���T�b�:��\ܫ�bJuu��J���?��,�5}t�jFgZ`��sM�.�T)��������%����*��	i�
�.G��� )�t�B�>�l5z�hu�7�ۻwo��+**vϘ1C��'�xB�?~ׯ��������}UUU�:t�V�(��ե�.��~�n\�#�<��w�ޭ[�h��&���2�nݺ�ɓ'c�4Q	㮻�ڱs�Ϊ�N:)o=u��7h�`�M�苲��*�e�.[�.�GH'U��{�0iҤ����_R��)S�^�M�Eux��e��0B:�2O���{�.C��!��XOF�A�:I	"���p��KH��J��؄Q��z�B
Q�| ��%���W�z�R����Y�|ѐz���Y}���꣏>R����2H�@H]f�2�8�u���v�ڙ�}�%�<XmݺU=��s�w�q]
)�#!d�.]]W^x��놄]�v�z�G�V�Ըq��QG�^x��e��B���i�K/�T�����A��۷O]r�%��/�T~�\���t���Ո#�OW<
�lРA�5����w�8VVѰaC�N@��~�ٳ'p��5�)s��o��w�q�S�N�A��j�*���͛�Jkڴ��ڵ��۷�j߾���Y�_|���O��_m:�e˖�[�n�NPM�4Q�w�>�^��>�o׬Y��NB�h6j�(p���-[���\-_����/]�T͙3G���ꢋ.2�@d��O=������_4�Ɯ��"��رc|B;���nܸQ�w�}���wV~�Ν�����J]{��U@�x����m۶9�۴i��+��R�w�y�����ZAg�n0}��P2l�ЦMu��V.�ݴ��%��c�=f��>}��jw,B���^{�HH,X���2�s'z�{�ܹ��o��u��O?�N<�D#]Q�CdB�v�ء�}�]Lf����ܹs�A:~��S�������M�PT)�L��d2/�\[)�`^ R>���X�u�$�xLӘyXca�����!Y��i7i>둹'N{c�!�裏Vݻw7� �o~b�Λ7/�^q���7�>��c�dM��̩+V��{oTD&��p�Gi��&�%RAgq����dr˚�E��A���M��z�Ӷm���i7R�	A2D1	��9%ߤ���E`�`�	y0A�z���~��8�a�ѣG,�8v^�\`*�Wz�e��ƍ��kת68�A�N>��LN�H�A�3����O7���t�/����Q�2!t(�d�g�6�"4�4�]u�U�;-��bd���:��À��h��g�}�t0�S�t�=���
c����%�/9r�i,��իW;E�y��j�ر&�V2$��sPx�LQ|#�nt:s+�$��|:F�-4���	&��S���^-^�X}��w�v��A 1n�c"#� ^(���=
�k2�Lz��!�}:���_�ިE�e�7a�N֭[�I���^*���'��_~Y���+�-@�� L慴���^��z��i��7�|c:J��@��̂*��6�h�4�:+�hQY\#j��H�O���*gDs�1���Ju���HS�9Rx.b���f��,�9���텶۴]��P�B{���
�͎W��F��c����:�"b��!��2߻n�:�Ns�i��uG��R6�ǀ�`����u�,J�{1V��Q���&� DA:�������!J:��Hf;��z�!��@9묳�IWZ�2'�!�=��}	���������kDU[]{>ȵ� RP_A��x���=�\cx�B�@��HG���~���Qo��e�:.�s�G�PP5?���!�ߑ"H"E�s�1j,컓@j������$*�1u��`LW�.�~H�`�`-B���{�Fj���6"Q�B ���B�/��s�s -i�ۤBs D`I��ȋ	I��/AE�r4N�K/�d��G��&Nd����[��ab�y6�'�)��6����o�B�Q�-�]�i�!�B-��H
uD�͚5˄?�LaJ����bM�I� R�,����bH��C�:��ʕxݥ��)� ��0��#�8�8If�$Ff"g
!���BA} E9p �����:�:$B�A#j�VO�%��Πa���ċg� ��1NBJ!) ?I�C��R�Ŀ0���rʼ"�C��v,�F�*5b, �H��&���̷�QW����IȚ�o�q�_J�9���E�Ro�~I"���G�U֣�JTmQW�+�b��������wBQX-�^A`��5V�K8q�%I��z2���ޞ�<Br��+$р�B����d1K�s!^}�	�X*@� !C֧Kv4b��}��wB��E=1�Ӹ�W��^�D]��-��	!aw���e�G��LrשuYJ)�I\�<�F"��ɖ��$���3L�6)�=fo`'����L{��`�#�@]�k Q`�[�oL1��!ue8���6��Ta��$����	��(��Rn$���L�X��@}�2d^e1����ӅT�FV�8��T�'���.�����|p	 ���A�~��Ǜ�H��,����Gbv����I�y���D�
�Z5a��R�B>��䄣$�q	(�o��sYargo	Y(�Fu�C~g�1����.s��d� F���D��Z
�= ���aU6�F"�0�X�bmE�����I,%k��bt Q�l�K*ܓ!�0Ŋr$��I�TTu�
I�n��R���|*1��9O|9���C�
D:���^�d04�D9D����)����i�g#��� a݆�"���$��dp��VV�;>I�L��<&�*�C<����wb0{I~�P|��,:2�B�F��0`�J���"�l�С�g�1V�D~�$E�q� D�� x��ā��4vQ�"!4Gk�����&S��b�/̅�M��5�'�q`�s��������&�ȩL򘛢�dz1���{�
���1��!�h.dp@Y�K̩���p:����ϟo<y�����	�>z�9���PK��'���x�^�O}q�`O�NY�lY�\lb�9с�Ҏ��E" ��;Q8́e�=%�|Q4B\'+D�	̉
8cC ���f�o�ϳ����>��9��~~��P�}�g��I�n]�^���:"���X*4�p�MFhTH��A�1�GZ8mG:6�t�#�ϧ��J�s-��B�S\W�TH��� I��ﺄ�&�
09r,'����h����9�.�!-�;U��H��ٹ�YS	S]"Mr-���	�Āi*�݄W��g߈b���|E�˒��� B���gΜyЙ���t"ǧr�����$���,B,2�$�߁Na~�_�A��A$�I�	���P[�:W����{ϼ!�49Ν$��w����`F�r$��?z�ĆI?~|A(�*ɣ�!r1_�ٶʲ��u�# dp���rڴiƌ���zğ���裏F��(FG�%����� :=�����ʳXv�G��B�t����� '.n���i�\�pD���	�����A$��oG�K	2R�]��D�*koG@�r4��8a@�P�D�#"�	8Y���eaOH.�ԽPp/�]T�z;�db؟�e���ӕb�f��hC�9��a��F���z�d!�3YaocNRX+�)$�:k*�B�� |"�X~��?���p!�a�r,�.+j��h�7R��(���}XK���9�F�����^��Ȇ��#��"�A����E��8��fڍ$��TNSu	�zo��S	���Z�U$�V.@�^
�Ը@3��x�i��_�~�°6�TM�y7!!L��Qy;*o4���*���h7&;15|�҃x��Hưa�bB'!���F�2k���mcƌ1VX�C �u�]�|�Ac�pN��`���k��RWa��I1(�Kv�!</��C��ϩ�U<s������:k���7�5��C�`�M.m�� 2述�r:	!zɼt����p^��u��\�D�9,��Y��]��K��,/u&`c}"I�v�!���NB`�;o���D����T��%����Bގ@粫
� �k7jU�z��qz0syh؃d���	����A$�#_�B���oA�D�vd^��z���,ƤҀ���gy�qP���2I��]���;��l���Ʈ���R������V���-��,*�f]��=�J��a�&O�4��@(��*I��[U�!���3���lP��2�����R��� 2@��UOJ28��2{�I�@2@�RO�8� ���܈�>J���wueeeϦM���[�ӷlٲa����U���4��iӦ�v~+��O�cǎ�V�ZV�sX:����aE	�ߞ�Kr�y�7��9�����׍��f͚[	�'�'�|���1��}(������{քx�xَ@n����Hk�\�"P���d�E�>p]�lՙ"��;�4?u壦���}��������,YRM��ɓ���!�~	���,W�"j��
�^���?�LԥY��%~�J��e�.CC��Q��]/����$h��g]f�Rp)q���ƒKtሉ���U�ž+��Ù�p.�������t>�.��d��=H��s���1����t�#2�|���xE,�Vx    IEND�B`�PK   <?XeX�^Q3 P /   images/a8051118-2cec-4f18-9b89-ac75f15be4ed.pngܼuXT��6��PAP@�F� DJZr������AR�A�F�T:E���k�ffߋ��~������o��������<�{��׊2$D4D�Ⱦ�T��˓ti����h�-���sY�����q ����K-G���4WSo�q�z�j������	����inc�h��΄���4qC���A����ܒ֦��2L�puy*c��,�YZ4�������߱�${}I�߷��$�?K)+_2��,�LR�qtKxK��+k�C����Y���R�JtF��^
Bl*�β��{�+��>��N)5X�_��zT"��5B���x�2ˆ��E�	��Y}~�����;�/�=���ύ�l��/�Y�zJӰ��0�r�|-��x�$"�A���P�p|����Ƈ�.fY��xJd��q>�#�g���J�>�K�6$lGȗK��S0�'G�xT}�3a�7/teȸo����\�b [߳1$w�#08}'�;�"h�������
�ʴ^�����i���0��oaot��R	{3��Re�2(BqrIs����:I ��w���s/�7ѝ�P�gG���K�\�,#�m��O)�$R�WF����%eLv}�U��o��������M��������T/��RB��N�cG�ы/JV�P�þ$�̲N{{�N
�1��S������|����(/-�.%����WVJ�wdoU��<Ҿ(0;v�X�xK>B^�\���ƪ��\bPyiC����Ph�]h�����ЊM�?)����Q����1-~�%wUO�jE��r�7]��Y�)c�+����֠$�S%"���K?z���WhsH�Ȍ�9F0+j��Z$�,,,,[�@�;f��V̟^eފ~� \��](]���ߟ3d��s_/�.��eQ1^&�\VX��Y=�ⓘ;jg�"�ѥckWP\��#��d�}]N�]NZ���_����0����H[ZZ���K����MCMݰ�w�4�r�j�+sƦ�����?d�f���φ.�`�w$��kZ�.g1�	��x���k�0���&�dfa8<<'h����B�D �݆�$Nz�y�AXZZ:M�T�ʧ��:�=��8J�5�����������d� i��Ҥl̙e>1!!��FX[[;-?�}||�wz�?8ȯ�JA���U��,ܼ��Y�.:;�`��ߺ�% i;5ES߹��4�{߶3�PӾ��?9y��ںl���BOPJJ���ZҊ�5�W�<��f�9�����������6rss�MVL�m%�!Ō\�Q�����.q��\\���M���������ݩ��v@>��i�@�n6�fm���5EPk���{Z�q�e�H�;��C�Bm�0�헒�O����T�gw������z�A�&ah�`��Rf�H{�x���Gܻ���?��fF����㠠2U�^e�h�=��Bғ�HfG�����j8��˹mٗ�&~�ȹ��eo�=���0�5k�h�S1�f����G��?�)���j7x8�/���Y[�	2�tqToll�x	�΁��� �Y�:	əB�.���i���`�I�EE�F�d�3�B� ���tK4�f�R	�1+���2>� �� ���/i ߞ`xFjݗ��������_�眱A111����Ff�7�Pt�|bbw����;���;S�)�K
8���~�F�֕�*++=�APp$l���8���ɉ�������4���:�ќ�?���mt}���Y���[��/9d��ʕ+��J��7d3(������R�e����:��bP�u���^j��#��vr*����qv�	l�����X=W�poe��co�À�ޠ��bU3S�5�>�w�AWaX�S%���YF���3˪`+:�j@�C@���Ahۡ�7�F�b
�6HĨ�j�фuU���N��eȠ�N0ӠE55u����'��l�F��|��,�E��lio��?�l9���|�=o0�*�.�ٖ ����[M!���Ҝ����N�ڌz��ps��G���J����c�ӸP#������_$����F`�!\2�]�i��L�9u�'l�ޠ?���W@�0ñ%Ӣ�$N�$�%)�?j��ϯ��1(�r	�ɔ<E˽� �ˉXLf�W\̅;lCHK���)7S^�����s/z(c�l3�P]1A�]�mMMOt�Ѳ]P����r *��&_�0P=_�����j����HW9Ө8u����=��ɉ�@�<_�8�� ��թ[�Z�����*@c��C�vͣ����M�bZ�9J��l�1�L�fI?D)y����%UX�H �e����򆄄����N�lW�:�IHI��GA9���`����bq�~2&��E*  (a�D�辋BĨm�8�L�/�_����eZ��Z~��J͓�Wp4�@{���\�(`n�� �36=m6�B��5�0L��O�����.� �肪>�,���UOsD��� �Ν;cK�=���ݶf�L�X��Y�t~${J�$V89۲�_�d~�w}�M�9���>�S�_�N�4���U܉̎����_bѷZ�H�����پ�{������틫{Dݜ [�&Fm���x�5�Gm],�����7w�θ�!j&D-O�Z,�]�f{8C�k���J3�E���/���ӥ��,��luK�Hڋu�?�^���2�6Y��W��蚼m�31!И��]�C�bD��	q�%��dA��I�L�Rb=��k'�����5>{e��O���������:�~�#@��ѿӘk3ezz�':L�By�#��HW��z�΃�c}�A^?%�ۤ��t�Jr}*7�<
T�(7��e=�S�?tTU���9��${��0N��|��Ò�|���s��͉#$����Κc������M�p���S��*,��C�z��ߥ�/��j!��i����Ǔ�C^9�j�WX����E��;~x��}��ߣ�{��*E���Pu[϶��Y�Rת��)DS����J������ۥG���/u����6?�t�_:^M{{��p���Wå��M�*I5�O�P3̹Ub֗?���IO�{w}> �,(�N|��φ�h*+Z�&&0}=
��� {�������a�'�ʱ����Bs�_ 
�Ԉ�V>�Q�x��_'U�@@�
@
_���^%`�i8�W�x����ʇu�fp*J5�*��W�p%���N<5�BKG6�2f� P��8���n;�3b��_o��o��z��j?Y>��VK��߷ ��iJM�������Y��{g�S�;���kr��mfD�d�+��
f ��s���O\ �n�#�NX������eB�<	�ңH{�8�A��paX	hﻙ�����_��D��m��c3�B,��'� ]�۸DǍL��h��*�C�ff� ���\�Wv�D�AQߵk"�yǢ*�
�f�E���a�% ��V�`h����T1�x��H2G�*�X��p_��ʪ.�S}��s��	@�p�nU���B�jQ]��߭?H�?�6:S�hi�]�$�Ik�<�X�
y	���i9j)��C_7��J߱6Wͮ0�j� ���������`���l�R�:�x��I�`OZ��߽U#ܙǉ�է�S��U�5�E��eM�ƀ[��x��o�`��{�穅���CM�~�=�^�PU�p�6��OD���v��wb}�	C��n�&<NG���B�ߵ��R�s���N�Z�R9���1��WQ220�(������|̖t����|��K����>�c��{�F�A֛��͍�?�R��~9�-�JH`%#�0�) ��]�9Dp��u�^0��::_�Hf٨�yV
"������m[��&�(�S�5$U=�ބ�q�����&���.��̑�=4C�:����������U�-���şHHH�Jc�"p�n[AH���D�udG�v�����[�A	����ٰ<�~5�<�g��D��(L\��KIz���\�m�W���m��Z7<������m.%0\�&���f�m7bC��q�����	&qf>�4� �)���ܘ��`�l�r��4��?��'�g�VRb�:t|l�ԙ��6fNHn~��fz�dD����-����5�T#u�o*��&�0!��ɮҙ*���Pb&�F>|�$�L��R�a=�����g�&+�y�㋇�
�^FN^�Kf��m��G!OA�2x}�.��i w!��Q�Po�?꾘�QM=V�_���Ӯhld��FP��Ã1��C܂pt����΀3��f���'�A���x�����8q��F��u�__ z�_/�P��U�,K2E�F��Ñ<�-c�ޓw�g�T�%."0�Uk����	��&=�(���|���
0��5
r,� G@�`�����~��cM�F�iU��`V=s&q%��'0ſ�����[dl�r����I�7c�X�r��lQ�F`~q�H��vG��H!�4���v�p��v/Td%g�u�[�Fc�7��O���*�e>��N�JD���~\1����=@4oUM�����0���࿁@�YSS�k�C�OR�Xi���I��}�˨�<e�4��$۠��*Z�J��|Vu�0�ƪ�gKX��o�V-$��y<\H
	p)������/�\�~�;a�_���C�4K�����������w=��W r�tʆk��-�g�W�nn�M:tqدW��A8u�L����Խ[n" lV������imp/p�A�#'�1BŜ��"ėt���'Vh=�$����=�շ���6�G� �If��������B����@:�!2����f�eSAP&��o��<J����+�s1+�s�4��]��"W-PǶ�IQ�����j�)�a�| {N���sV��s�a4C$ڟ>�=^��h]R�2�`�1�q��l�*3e������>�����Nv��zPu�0&��R.�hӝ�d8��o�?;��b����qۏ���f�Fo�ܘ'k�FN>+���+�#�>�!6uE5	n�c����`Y7����P����q8�&q��&�ڀRa���q��%FH�궂S����$y�7-����r_���>۟����f��x��^��`����	+�Գ5S�X=�;�!+��<��\2ˋ�
Y�З^P�#;$��=��XBC�\]���mQ�TH/��:��{q���oܐ�YV�V ��YQt�";�E�
�3�H��O��2t%�2Қ
ʹG }�_�$v���[U�o�1�a���q{8S�YZ2�~�:�gY6fU���_�SmmmkJ%�y�	"�c_Pƛ$�:�����=��|0�oS�w��|�ag���uHI�2Q�zz
�����Y�_�,�l�6�Ku(��0��P�7��1:�JdlR��^�h�2\L����E�2@M���V��v��q˰��f�ɛ#H�7[�ŤM�j���Hdp(�� P�B|/�F�����G�U�q[a���P���/6��iC m	�� V}�#S��5�(����|��v��	K�oP���f9�`���,`�}�3���Ǉc�:��]O��Om2.���\(��mbuoU�\>r��E.����9H]�{��d���-��wl�w���|'��z0��,U�5%w./�' �y��ْ8JQ%�u�7F����x�Iv� ��2�{p�H�y�N1�Q���r���Hљ�MǕF�w��)V���@x����O���D��dV���eq� �P�FN(#�B�=��x���?��R�~�uɷ�<NS{��}��{S�5��h��;�.慉̲��mt�bᭂ�
�ҡj�#q�~�T��٩��>{�m(�s�g�%u�6���m«�ЏC (���h�{-�e�ݙ��m�^���:����?/U�x���L���^v�V�ԨWʧ-ʧ�R`�A��<�[��-�>hF���Μ���~>Z���j�V������&7PNKXl�C��¸���z��tm��2>B�J��H%��XyWn�H�>�%Pг'3x
"?�|b�\�K�t�666B���oՎ4ج�XVP��>R��Z�S�9A�� �_*�L��ܳSo�L(as�����zl[���xa�KA����xvws֭�B��h�74xw����~�/�w2B)]2��:��_r�>�L�Lh��Y\e)Ў������68���L �>P�<"""�YYYB�K阦��wg���ZF
qX\�iMQhJf���75o3�Xm�Ԧ����W�
�nm���i`�F9_
ؔͽ+k���~��n�%%x|@�mi��h�������5_��ĹS��F�d9���?�v!q��1˖�t�G0!���k�2�o�C\Sy�ُ�\L;�Gf�?��\p}�Ԛ�ڊ�z�߸���m 4|}�-���
�=���<
u��:u��#q��qr��g̪?��>�Yh+Uk�=䬙���;��!$��*󖷷7�V�IlW���S�&�?����9��P���>����F��@ߖ/m��sR)����,6�����z��<��/�r�Y(u�_e�\�B���6]���L%1�u�:=̲���A���Wv��
l��W+���"��{�ng�H��8��~�r���{��f�Л��d��jnmRn��qv�k+S����3S�b�pϢp#�@�6�4H^qgb�vr��@ir��< l}vK����_��������H�G�]�4l8�/ě�z�ZTд�q��p�	�P��Ձ���6��K_���aTú�hλ�þ;6��{n亲Ce*Y�"o��"�|�B�?�����|�2���?$8X��9� :�4L�[uE�7�{:O�z�� ��\ڰR{�V� >�J���4�[���J;a�l.��O���������"`W��b�)ٳ@f��+�9�\��n��Y>h���F�}��~V��dV��� m?E��Ρ���^�A�Q��уuacY[�ŁG�ɴ0�5����xS/�=s2���/�tz��W�c>m}�g�j7�(
WU (1,bF�+ ���$@߄ۍy�c���e�ض�u�\�R+<{��8�� ��$.3��)ꯞ�Qn�7�<&Tٸ-�`�<҉�������R@�MM��Nt�豢���Z_��	��8��t�ڄʄ0��7pѻυ�INLW_o��m^L"\�V/�:i�-Ӷ_�>BCq�{Ѿps���d�[O�Y�=x�V&�S�I��Qӻt�0q�iS9`��U.'���d���*�л
��\%�G����٨f:V:J�)}�ti� r=�j��Pc�îN�Z����?(	�9z?3XG�{�c`����GԴݸ'�Q�,�p �o���@ wȢd�
����wj6��<��]�:XP���(�n{d��l_{WMNF6���Ը9��
Z��j����!�>�[QU��[��}7�ϩ��BI��9�-����������@�������KJ�����e�x<����DkC:��?�V������ ���3��ס����e|�\�4�3EӅ�5�MO�FPA��|Xұ*�O��\ǩ'Ƅ9�R<Vr���Ubu.>M����V=����)1�h_ܡ����5��s#ӏc����j8c��U(����+�R��p��S���E���I��9sn5�Lg⥣�)gu��=�ӿ����8f��x#RI�ķG������%�	$�n��2������B��;��޹JФ���v:��� #��ӳd� �vHQ�ޞ�T��o�t�F"Ľzur��7R1`�ÍW����b7�g�t�=�Z����=����VT�BU�ש{7s��|(9�db�US��2p� ��mܞoG.��
rsߜ9l��D�^��)D>��� ,-��)��-k��n�ii�)~�{�G��	 �q����J$��ݟ#37[؋�W��T'���q���l�Ƿ����'Pa�r�	�	�����`wEm��O`���(v�V6�B
��ON��]-?�m	��Iݶv҃�1R��Pۀ�:!T���;�}$#R6t��0�
FYhqUU�����d	���Q�6�y%]����)·��ч�7č����V/$X��A?�XD��|S�N�?�* �z�%�&��k9�n���3<\��mA	x^8��^DPq�؜&fo��ӝ�
?x�:�\3P:����nn���?4߅�?���͍zn
��TZ�;yu����9�͎)(�D����H�V�v�.�s��W�5ώ� b��6neQ����? F��嘇`Ӯ% fc����ۿ^lu㰩����@��} ]!WR�(����$6�eSw���_�P�Lp�0L������@bHJJJ�cܺ�X5s� x�>6갍!E�c��K5��f�>u�ڗ}{4:bц��/�I0��N5/�Yv���.�R��g"�^k��9W,����1˙��
kk��Y���Q"�F���kڃ�E8H�������p���W@��&��I%�.� j��;~��Mݮ��٫,��ۣ����!af��X�>�X%��9��p<�80YA��JЃg3W�'��M��b�?3��wV"�GK���˿3퇵L[����8� ���)�<��,Z&[f��n}̟���/N��	u߂�'������63~�hKHG�2���S/Y`b�உ�/$��`Ad���G���_��d�Dk[�#��wu���/��8-?�r��n�ќ�q�Tl��U �b4@�:�������K��������&�^|�����@�ok�0#�����јu�i�6(�Q�;�'��Cx[��V� �������,�����0| �V�04zw~����&T%��tˮy�I��0{1���WF�+�%���m&��s�W]��b�7_v���a�Me8�^��*VYc����x�r����4��C�)y�+i�Z�]?��6z��u��xn��M���r�d�R#�FN��/���������-5���4�WA|	w6���,����5�W��כ�����������]
��	�W�,N�lC�Q��y8����?���W��/��|@��B�_�~]Z]�����$9�~Ҭ�����Y�4��B~2�[~�i��ځ0c�|�5�u2�,R"��~ �ב�q�����.)LQ]���&�������Ęo��m5�)�r1��*/6=�i ����{a��כ�;=��3c�)nx�0W��?2�g�,��%��g�w⟷t�5_�^�[M����+�\��c jD��P�k�<5`�&q�*d�е��?1!ZD��{�^�m�������K��L�O �[C�}}{���y`
�c�8>�|��ў�\	�[jg�"uF��+	�qN��m.����ړ�:̿��]�J�����we�SSt����aͲ?퉅��O������`�y�����n̈��T<����cȧZ����kJ[9�ɸv�{�	z���q,3\��¶���~)��xӔ;/^�P�&���A�ҳ�YJ1n����4޽��)1��u�:5��0��fC�Q-�_�^�
��ik�/J�ݩ�mm������4�M����ύ����}����jg�fm��N�A��e�߀���<	�,��U$W��+q�v�إ�%����|(G����Ϩ19�ӵ�T�>��x�t���b���>�i�H%�Kj�T1���mWL�n���V��-�DpO���&��J0�m��X���]�f2��U\`r��vW�[��+JhE��!��a�-��J%���Q]@I-�����4���]\�.��Q��g�#�PLBB�HW������>g��wB#����]��N�l��I����vi���O���T��M!/Qa�Чò��I�"��|{��� o�T[�jQ_���z� NW]���b�=i3����O�++��{�i{3ƀ�<����:޳��[tln�]�|'�/���Y㦂�?��H��a�,˛	��ZS#���ɔ�VS���ޡG�G�YCz��yE����!n�S��.cx7��ǋ7]k�-W�gg���?���I�=�	���F���f�6�+���M�y8�d����0x;
8`5&�w)v��6���AF����c�zW�;|��NɧZ�43��.����htJEMG���aQ,)n����� ���ݕ�<9���r�??lkjj�2�E�;v<t���|�:M�]a�}��k�dejj<�j�����星�d��3�QFb��HJJ��EK�U�_G��S�u�j�>#�Z���]��?lC�s�s�E�kބ��Ol��������)zS��kj�RZ�a�z���ԁ+�P��#��N�O�K�� Ԉ���=��y��n���RR�9��8nKU	F�������ό�a�������"�gn�t.KQ1��E�+y�+y��wP^Q!Z�@��#�Ȉ���/�I���2�}����ws�
%x�88���oS��2����@b�	G|��#�#������C��u%q���q�� ���/?��}#�K��W�I�`�j5�k�M��,|�p��:�!33HKK���j]5u��KB/OS� ��?z�#<X#�v�����[�\�wһb2�5�
1��/�6:�Z�7�ٲ�n�t0��x�X��{��4���D�%��H�:��0qa���7û2G٠�?�p���A78\ [B�ҵ����-��l��m�{�T|�W�0�=�~p+=3�Dwնao>��O�������qBLzUؙjt `@4���&1�$�����Ӓ��e:�{m~�b0�XR�~�@P_v]����h[��X[�h���x�"��E��������r�K��W'���[��+�w��˿7PI���U�<>��'���zJ����|z���ǝ��$E�R�qK<V�VG��|)�_S�V��Yd��7�>q6��ޒ�Z1LQ�Q�HeHG0�ok
6n�P��%��Uc��L|�q <����O�av
��蟄�t.XoA���'.�ʒU�Y�}{�߸_A�#����d��v���<r;�����R�(��p3�F��_������D/+�8��e -�i�����09�#sp�r��X�4�{�2ix:���1
{�Μ�HG ���G�M��p2���0�iYՌ�I��{I0�/��|���/E��,�U��~���v�������n"ѵ��q#O�	"��N���/ �|@��h}}���h�L~��|4�s���ac;ZLe@�X	V?�}K����)��|�������8>�FP);�P�1��z�9y{˂2�*hJtv �$��녪�E�B�.���on*`N闏W����$<>0����[U��� �<j|�U�S�͓  @�3x�#ߞ�)��g��/�K���쪇-���?��4"&O (��朙����cύ��k�r4����"?�bBC�0NlW��Xߋ&V�;::�lgtX��KmEt�6�j �q�A��cb�M,�!E��%ymw�X��@�� ��Tu&��g�������~\)�w2���Q=����`��A�,��SO��c9�r�|��X	lT�����z�?��M%����� �:9;K�ȴU� �w��xS��,��ɑX����زpz�*i\'8����f��^���@=§&��>�i�2޿A4,���@׀Պ��,4Ϣ�c���&P�)���_1��gZ�W9�z4��&%��]�2��/���l����]���~*������5�����.���1}'{+���E5�։7�Opz\�aɛ^	Bj2���Sa��"���B���3^������_�R�\���E�'J��D���j�-�p��b�^Wy����>ʊ]�'X4RS�=S%W�ܲ/���/�_2�W�nU�#��AxC�Mx~q�!LD�JA_�������FrB��l�a�"�9����<�|���� ���P�ܚ#�KC_��pA��A�V�{+C���u��W\�����N�p`��C\�Q��!�xN9wڵ߃b����Do,t�í"����z�>Xm;���I^nn������p������E���,Zcw!v���o�?�D�%�Qg�L�,5�B�l4��IB�.���.���Ne��7=�As��9��"cZ�I�/��@�����)���Щa��hO�I�d��dy�������j�Nciz�������fS�:���<*��(�rn����{n�Ƽ����2a���_,�N���:�eX���t;�gWAl~Ğ6G?�?(�֮�S�^�m��=r��Iti��;F�1 B��gD$u�f��'�Bb�꧰.��L�=�_�i��AO+Y'�N	9����g��(\ٕ��
�\(��O6"�=3�%���~�1o�F���`���9��D��R��@e��-� ~�-�D3S�w4TX��:|b�O١m���@���+JfN�.��3�&��|�)�C��������yc<Xj~q�v�'�U�Қ��UV��N���"�2J�{Q?�~[�/[=�˧ڽ���-��Bq2^�^]׬f�=:���Ǽ��=�w\��ݭ>�WOj��e��|Q��l�@�l ��\���<Z�9*m�-ٱd�8��X~6�Ƣ�ѳ��0=u4� ���ݎ�ŉ���5lo���t�z�h��W�4R�F,$�)���y���ٰ�"~�; <� A_޸5L�֊���U?G���`��1��T�]|�y�?���=�C��S8����}�ɕ�K�|��)?�b��{�rb�{G�yH���C)����y���a�4f�$#�S��KC���p�^D�mS����e//s�:�ܩ��5�:ݦ*��t,��t��k̟��p~��Z-��h�x
�����)�f��X������d7���k�ع�tF���;�^���`h�9s��\(f)����;Q V�$N�%�4��_�E[�q_W��]L��/���L\p{�5n/�^ �����;�7��Eڛ �̎��=�NQw�}׻2��n���ӭ�5Rz��v-�k���/���n�t�)!���k�E�`=�K�t�2�՝�d<���Yt�pW�]��^ER^�;n��K�S:�ήY4��T<꼟^��a�����i�1Buz�B�)^۲@Ț����M�Z}8�Yx��ɤ"���26Snp�U���Ψ�w1w9�t5q偂t���ܿ���c�ާ��J�z��n�s8Qi_u�S���P_��q
��^��Y���A�a�
f�|��-}s;H�g���:��R]Ԓ��~�����V�+6\{�\2����"�"�u�ٺ��9�_Q71�������;Jl��w})���Y6B�re��(NR3�u�AL�D�����V,�56�t'�-�k{��1�@�,�Q>j���ӣ"+�6:ץƓG.p���6L����	��/Sa���p�N
�����T�LP�k��-����	��Q RG��[����<���í]>��7��$O&���&z�.����h�>�Ҋވ����!<wshxx�ݰ�]��Œ���z���VQǏ6G~��YՕ�ke���O�&�5���=�0{��(v��C�ް�������-<[=u��@��S��M���+��4j���,֞wQ��������o��:j��o��h���v�?R�md���ԝ�Ezg���3�;`��x9����2p��ꢼ�_�M"��VNC�������db�r��C�:�{������g|�CѺ�ݢ�J�YMT�9d̴?�<*,���3��Ek��?�e��ssr^�Ѩa����4iߖ[\l����HE���;vz�K��j&W1z��?3p��[�6ޕi���L��̶"4��=�����trZs�ӱP��FR�Uا�TW�,���Z�ƄN���G/����1�k���|��Q���¦Qv��3��ț[D�X�CN-��@ܺO,q\,������ɂ �F�|�� 	�t����ٻ,��B�l0�R7�UJ�x��8lfѕ�
�:Ql�%�FZ��O	;Y+�Ш��v�8��X]������gĔs��}� I�t~ecC 
Nt��VL^~>e���2�����"曗���x02�nB��X'�>��{.�m+�ώ���8'���*��'���[&�(JH}�Տ(7ZX���ω������{�InV����W���������ԼH�哖4$��;I3�.5�7Yo��`�׳ 2�+]\����)�$� �
u�{
��k�}���QG���q0� s��͛���R�Ò�2�^����*�pC�l�$:��mӰ��GR��E���][�Ṿ^!=�ᾆ�� �Փ���������D�����N���J�#FqM^�2'�K?R�U&� �������ͥ�3���U��%�z���YIg����z��I� D|��9�!�79�h�����V�!|��k`z�0�-}|\[+��p�������6�I�5�{�Зϯ��FŌZs����қr��[7�7��䢖��<���{5n߷�'g�!�#�/S�~yb9|���7����7�ḯ��� �Tἆ���'�h�?���Ү����J�IP��8D6�������_� D�&�/�7&ne��"^Q�zw�A�����å���n22\[�=0Sܛ��z<1S�vn|�������{3~�﫫�W�<eI���
��S�_a{��	U�@D��D?f����.�����ܟ�,�G	?�R�ם ��g�iiV�g5����n��kh�������Ό���F~g
=o{���|C����c����x�3�
|���gˆ��ն�~��4b���sŅ�O5,G���e}���+7 bl��b@�t
�ݥj���y�U�W�1r%2�m�٬���u�,!�ت9�ea��7�i	�
�I�����X������s��>onf���S�6:���;O�;<�7U�׬�]�ߙo6<���71>Z��>�������ί��p��J�r��]L�2Sܨ�Z=_M=��f��X��w6S�w�D�zΫ�<�L7B�D���i�/泌�E
�}0[:;g����wwR�\���0�~�ȫCI���.�u��Wf�ǅ#��^*�^�~=�q��dR�0}.�/.�����_6��|�~�-�0�Щ���� ��X5�p8���D��L�,�1*������^;�-��������Y��+���k�}͚q�����p�_���uRhac�_#Nu�����.F/UT�괳�#��X�/��!8�`�Qs���X�h��|�~���?�4,utt���j�J՜���{RUD�� 8��e�=����պk4=,�mn�xn�~b���h�+I�c���*S�H��8�e���_�.�#���B��	�vr�����c�D����'��.�;wמyJ_3����
n�0��H���tA�?f�a32�w<ni[GI}&d��/��mD)r��*�xwO�=ڃ�H��1rHz`�6 �m"����06��e�l71?�D��x���I���M::" ��8S�=�;2j9�QΉ�'�׸bc�߿u����ק����坧8�yX��֖���*{�l������ݴ��!"�nۢ�<$�r�&�l�{8�E�E���q߱���0|�����R��R��x�j.�9m˂`���p=͎뭋PP���u����ml�l��w@M�a2����I:��o����������6�$O���}!f���Q���f�ZV����i���^;�����3�������ć��`�W*!���%���$ϡ�:��V��;Y�� ��:6'�A6�7�������<�� �E=rDmU�j���������1�C?�b}��Z)� ��&����\�9����6@��h�9҇~u͛x<N���	��?���!�G�e�"r���@fp��=�MYt��5ݎ�'f�ƭ��p�9!�H��_T䆸��F�C#<t�������*�;i���E<�s�{��c���Lf#y
�KR�?6�VL���(���GLb�3B�,�Z�R/���<�������i�U�s���� Ex�jvu��[ی�U���c?E1��I�IȱmM��$d0��\1>w�x>�7^�qtuZ�2�-C�n�y��EYs�H��~�H����Z�v���>�õ���,W�Ԕ���X2�-�q¤V�Q����X��,��+3���~\��������>�����iRL�`
���c�we���K;�S�9_�F��槥1�W|�|.�X�Q4���f{_��!.�v��ɣ$r�5+�i�ٱ���|�-��ȉ��!��?�a�	��WV
<���`�K���&�{�1�����/�Z����t����V�w��G�U�8�S�\�ޟ�b��B��9�yp�r�D����:�]Y��'���	d~+��9�L:Q '(j�D
O3�/F�}�|<>��Q�\X���)Y=f��ҿ�*W���"���ى��܆��EX�>���3�������5��->���iJ�7U%��u^��ع���υ����;2Q���_�oω��睝�D~�ډ��[�{K��NnmTĮ���ky��_��N�.U�����J����2p}�(PF�S��u��wY.|&�������Bt������ڞ�C�25�J�1�k洔R�L/��z�=1�Ʋ�l�Qi�c�ޥ���m(�LXs�ٿ|Vy��c9 ~-��;VL��|���{�
�(�$4p	���؛rZfe�WN*��mp�91�
N���1���Hvv���Q�Ī"���uuC���蹡�B�X�5QsG@�MMM��45���щV[�� Ԫ���z�>��,���=�{#??�2̒��{�V�Cێ�t��"Y'y�)6���f1A�%�H�lšV��!=��`�� ��
W��]]]�3k�'@�j�Hy�$k��%$&VXOT��++����$���X��KE�G�F"}P-@f���`�S��ߩ����v����"D��y�����%�O�z��-����oQ=>�3����p^ը��
;�t��v���R32J�ݪ��BB+�z;h}����}�����v���*�ja�3�Xq=x�>-"��ǔS��d���F�pbdE.		��8*e��uͫ =�E������R��������[��?岖#ES�[�Ï�Ó���/�r=yg��A��/n�~FH�1�\��J:�.Q�$:`�Oq�IeeVJ����֮J�1����[1u�)б�ΐ����R�N��v��BW�D�f�j?�u��D��Qkp���,������\�zk���	O[\�{���3��YB�//��ūf���U�tE0K�+"��ttt��b�=Iª


�S�O���_i��)dS�3ɱJY��$琕��8F*�:8Vv���	���-�ؒy̌��~����_��?r��������~��*)������_�B��O���<�i�)E����`��3CL������,��o4�i������?v5NN��L�م}�8�h�ř�]���
�Jcӗ�w���T���+�����h~b���)0��a�g�L�&as5�1�Ǐ�x�Jlqsnj��DEs
#�j���.+M@ �G3���������[?BJ0��]ؑ���+#��*	��o�q2� �%���,����h�z�G�ut��oJ�![�G+��u	����������cK|�BN�A��HX�m'��&HɈ�)�h+p%��a�ӥ3����Hu�V��Dǚ�K� 5���6?�~I=�)7%�^)z��� 7Eq�}��t�vss�v���g�\� q&�ۀH��Ҍ����7S2ҽ6u���d��lB�m-b���>�������7��'=rڏz��x��M����y�G��iȀ�z�3��!�=��m��+���t�o��?{�_��J��jj��8�������cg?7Jb���=1H�P�p�s��3R�M�']+�� (wEb�p��G��Zߝ���l���^��� (t�6�prP��ѸW������}�p�(4�O�|��"m|b����ܲ2���r˞,�.��FF��x��ZR˽��59	il\1������{��q<��hm�y�~�U~�����+��o�+�;%��i �PU�hT���Ff�p���:4�6R�m�&1���=��b��J�v��ž�hYY�D�I	��q�R^�خ��_��S��&����w�>&&u&�Ng{�S9ޕuΛ�+�%��$�ŒN������K�}�U�2�}�iW�����Fw=@�����ϕ��9Ǵs��7����O�RZͯq�*��D)��`�44O�&בxdj������w�^A�|�xA��1z��u��g��0Ѝj�[Ю��6��~�3;z2��$�!��������K7�g��"++�����H�r�s�;0X����6a�{��F�C��49,�_yͫ�h�(�r]'�������_R��������T��*�����]���ž���*���3���S��0]����"^q�)�y���IA�I����W�LV'���-*q��&4�.� ���8r�W����^0
��'_/\��x�<����ǅ��س)
}���ZSY�يk��y��Kv�\� n�Ȯ4a���f*�=�}-r�s�I�$'/��Hٴ����1B�ܬq���(Sm41w@:�h���9 J{^@�[b�CCh�t����g'����.��&1K����?1���&�;g���ҍ�^���諫��1��x�F�4,�N$�>�f4�5R`��䇵�}�Z-E`�婎-�V[�7�َ6��'|t��sm΂xVWU�}������mU/���}�v�zAF{�,W-4&L���,3ROTL�eM?���5)��lݟx��N�6���ғR��B[{��m�EP�D$6_E>r���6�N{U�3ZR�� �Z�ՁgN$��u�-��g\�y�c�{u
b�lt���Z�T�\�$��Wu���C�K�� 3����I��a�섕y��QP�����4�y!���'#��L�W�j��s#�s"j�0���͕����ꑂ��Nj�qc*L�#�r*
\��.���	_N�A�F�+~3y6ĩ�9�Yڧ
��祥=����O(�䰯��!Y��rU���N<�["2g��|�>����֝ �ݧ�\�wg}��S@�Hn�P��7�D��=��Y�/���|\>L�gk�Kn�lJ���o��ҟR��-2��V\RRbck+�D���,2�-��L�k3��xKSu��r��.�t�BR�r^�O�1F��@���Q��c��[Hs@s�D�H�<���\��5͔���z̰���f�[�����C]�H�>|H�v�o$9ǔߛ�z��x&��ȨmRk�b�,�ݤ�3/��W�>	�R �u;�>�F��V�w"h�BH���.���Z���}�`��kc������AQ���4���>��R�vI�}�����E�J[����ą��>����r�n`�����J5�t�:����H�� �('c2��b��DԽ�p�����EB�>Q[�'��w<�I��w>����)wA����P �\���#��ge���$��Y)B����5@jd��Ƴ�D� P\.��'�s'x��Y�6�)m5��bL�F�=?\����o{�����'D �kIOI�� F�Ywҿ���:����W��W� �<��2��-�;
��Z*��nw~�ސ��wn\
�����=�K�>Є`Zo =�ҝ�j��%��x)���w�k�9�O*����@�c�)*�r�����H�����䗖/:E��P�V��?��k6qsy�imnT�o��j)�f�7(��f���[��o �#� ?�|��k�u����F7��{��S���L����z�Eϰ�.laa1����#u�T��!s����l��O3��]0/]\V��#�t������n��o��H64.X�B�*�B���$��U^����O�)	xNZv���c`��f���s�A�k��&l�%J����������;]�C �?(nw�c~.W�%�\ް�t�iqG�*�fl�]��}��s�{w��dd�j8T�±f��"��pw���w3����l�֚5�	�����ø�9<���e3�����X�=>�y�ʤ����UxBބMsK4[J(S������ͩW:P�e��F(���:��u�h����;>�X6&��3��4�C��F�%j��<i�Eŏhu��_��o,���Շ����JQtj$mD� ��[b�T|5��N7�!3�O<�����x{�Rv���(h��V�S?�-���1M{��	s <�RY�۵� �wL���u���d{��y��^��I��󅀷��ɋ�+��	w�T���<=�ő���(sak��C>;ukN	c�[T�\/G���`����4�}�S����4R�7��$��w�R72��1N��=:ʷ��:���W^{n�YTC���^�ύ����(���u�Zu��~����rj�R����U��-�o7X���U`��ҟtj/�`���+��{���3_$[\[Ӈ����Hx�K�_ӹX�W�9y��w0�e����x�!���Ա�9�6�5F(?J�_]�T�e#̨���?�(�~�JI)��N30���@���js�F�l��i�,�6��<!�r�ÈJ:u��ת�������^�H@D��D��)�����,(J�����X�gгrm����VE }�q;yp]i�{8+���ϾG��,nTY�n��ƃ��=�w����Rf�]<���¤2u�m�^��`\�2����+W2E�%�Y�QD�ST�;�*��V��O	���U�p��Iy�^��6�Y�Pj�l�W���!���Bf-��ʱ��G�4I��?��ܪdV�=^RSz^�]Q&�[Yko� ��D�sǋ�X��n�����;ݨ��}�D�Dy���?��T=��w�O�5�Z�Δ`��J�R��HF-��{�nDg�O�ц{����G$p�2,�!��f@�58 ���ۊXrN�s҇�V�@Hz�����e[>�e6�Ċa�me��G��T-�����6�X_Y�9^C��ܑ�i�.����1��G�Jk��ʷ��H�.+iƅ��˼�"�ҫb[��Íb��W����E<�|U��J�ޝEk��T����./?uw�x��� d?C܃'����t%߿�gg8�^�Z� ��.�8�� ��"~�=��BBT�}����|���
��Tⶔ��<�v$��4�;A�;F�Eؔ


��ZH\M���u;v6{�&7�3W��#�O40��o+RsX�j�z�h�E���h�*йsp��mpW_�f9���B�.%�Ig��
�	g����F<�
���}�q{zn�����Ts�,3S@�m�[�"��2���_���B���δ6�|��=�D���3I��`�e��6Ov�aO�9q���� gu���6�,����cb���p:����+>'{ɞ��bL7Xd���@����i#n���%z׳��������ӱ��qVj���RW��7��҉�V���|Ǧ�ig+�^$qA�����,G7���*�Mt�yG�2_�J�9K�(]�Ý�ҡ�>�Ƃ=n�q�)������zc eT�� ��^��W��[J��Ð�+�~�Y��J��;�~=8�w�М�1���;���~�>��S7D���v�g'���h��{a��������a��_6I��u&G=jRD1�����x1G�ɡ�7E���s�"Ld��[�Ȍ�m��>�S��TM	����=\*�8���S��sI7��YQ�J����
�`S��iE��p�¸F�����j�$��="#,�8�^L��	XG����}#��������@�Z���9T"`�:\�?�|�ɉ��x�����>!ynS��B���G.�.�z���%%�>��Hŋ�#����-�yV]�\��yUU����M/�q���6�����>��Sh�0���|/\b�`�'��
�{�"�wO�;�OCr��I�/˧��+������)�X[GNS5�\��5�q}x+
Ͳ�ivC*��j�X���NF�G�?�B#-y��ؕ��:�o�f:���|L��axކ�nVi�G`�"��	_���Qb����<9:$��l^��4�C�p�����`�}BxXŏ]�z��L@�5��x�f#�.xV�5\�ah�L1�̘��\�v�V�t�3~C�@py>��y��4}w��V�?SV�� ��s��@��U�p�&�jE��k-��o��]�[?n ���3�U��RY�ۧcm.�M�6ֹBLf��eI��{<��-��xC��AT�w<��١��e�CN�<+�8V��V�S��Nr����b������E ��e��qս�b�gN|���~�����f~�!���Ꙑ��}ѭ��{��G��r���� }�;ו��R؄�����ɭ�Ï����	Z�j�^��O��?��EtӾQ�`S[�PD����|t�o_��(�Q�~�`5�G��4 b���(�#�Krz,oR$9��Al�����%�]�Ql��{�Yݷ�l�(�L-.www�SeX7L����,Z\4}'�u=IP�z��QΌ�e���U*�:VI��!���mlM'���5b �*�J =��~��>4~#[MeD�pK/�w�: NQ��[ޠU%O�:����U��y���<mp���-�OȤ�H;��~m����Q���Y��������Y>�8b�����P��s>K��Jb�.�k��Ϲs&�v����_�;o����Zců�:Di��[���.�bٻ��1Y����?�N�ݛ�yj����y�9�bVcSV�����-[���B(�����E	�{�!tI��}��˶h�O��(yk������zn>q^�"����?7�n�Hm��E0ZL�eփ\��6C�U?�6��Ye|(�y���O���$HKNNd�f0�؟T3�:\����|��a�E��9dNZ>�v-�(,��V�{/�2,��Sγ��i��ï�T�+��K]ҒF{��м�u�>�8�Re������I!�2�\A�ǋ�$ �v��f��ȶ�����g��q��\y��a _�w	Q��[=��U-�WJ)����Q���GN�ݘ�h�j:�H�FeX�q�1|����C�o񟆏33�yb�)Û�k��q5�ZO:��NL����� �th�� 7ǿog�90���h��f�r��|�'��DD����=�����e5��=,*�-�~�� m���^Hl~�	�1����Ev�$��#��kk^ù~�5��ت$�S)dRB�㑾>s�b	]���dTZ��	:�N6\��ڢ��I�G���AM��]Wm�<�K�s ��2 r<� �c���n�7?ʼT��c�M�ӿ��[:�q�7���L�٘�8��g�K���J�����
�X۸�S{ԏ[H����PYA(�=d��ؗ0�e7�(E�������v4�VZ�O�u)[/<*��|g�5���V�^1�q���g�� `�sAѰ�כ�kR��d���1=}H>oK�P�ۛ��ss�U9���_�KG�'v]��ܕ�QRW,�����DP �~i��]+�X�Li��`c����/涩(<��͌�"����ޥ� ����>*�؃($��?��E��H�6�*J�m��i�W�}.�+��K��Xq�*�Ap�x�,�e��th���&�Z�6�꯽�n ��Z*m�Vs��qsТ�3&|���d�'�@�����W��]]���םdƟ���;�����Ԅws�~��W�<��XF/=9g�ԖQT��ϫ$8�I�4�����7��<��ʭ�p���B�]�N�ə���0&#11��svJ׫�bf��vV�1�~t��%�G��9�{g}C��S�vVKQ���H"�{Z�=�`�.������#^)G�,�(5f��M�� �M����C�ҧфӻUlR+��5���=[�c��-%$2��s�>,�s[�� ��Ɨ.��������^��&��]ثA�^���ԩ��ݥ��m�,P����W����7 �5?Zz���ֺ�y+-��P͝||����Z��U�fΣ�G�55�M�I���c�M�$���x�w�R&�FY˵�%�n [$���"c�����1T��9XF��x�;r��-�����ک` ��q���?~i��.����6K$:��S�����ƞ��g?�@�\L͛I�ŷ���mk�X�k�~������H�V�_(:lXN�ם�&���U-��%RJ@ KZ2;����H�7��n�t�O�6+�X{����0��p#x��㲫>kmӶ'����̪��ri(������y���/��*'��_��Ns���u#_d�	�&��!��h�&j�[���2��X������.��jj@�&i�J�o�4���⦃�9���ҙ�dY�<���}�������u�x�M#N���h��Ĥ�il��U���v��l���4S�ˡ���8SP]�9�tS�����T�)�l���)��,�WĲw*�-g\̆\Y��v�	�S�|�걒�apB��"#6�0���`!ya���&��^9�o9w��:�3��o[�)��VPvjl�
�m�;e�]~t��~�
�I�&٦4�).��Δ�����8ǘ�0�s� 5E{*ɼK÷�k�qG�+'�j�Y:X���ouɴ!(�~Fj�>񾷠ڇ���y[��g������~wδ�u�HXѪ���;:܎16�h7�� g��x.��K.�Aұ&g�R���1
�2YH�
W06[��t�����yLIG��\5Β�����}E����􌥌�ؗc�HbJc�p[��!;��8���);9���3��6F���&	O0M.�ćVVU��$z���s��8��᰻��\�r�@^�s���gZ\PU�tGP	&�������� �7CY�h?�Y�q�0�$|��.�3��2�|#,
��;���#+<�	W)�[Be.3%C��%�;('��=H6��|�S׷�z�gjbCB�ӞL���Ís~E���`i����>r�����#V�K�{�\�<�p�v]�0�\B��~�rIٝ�ķ�F�-�o����у��¥��q+ޡdڧ:��	����#�U����1�k3�+����o^�yƍ�����u#�O2Ϟ�%.]��lr^�8y2%s'7��i���l-.�s��>a�9{o���$$|D9�e�آ��Ҍ� ��
Rqƨ�%��!�?:ZHݭ��!�;��1D��aIפ�,�!ޠ�g�]�N=e g\��Tr7���3�W�����W���n�+�����sO¦��R|���Oa����;�Q}=� �}����] ����z��!ʿ(WFR��,�9��ׇDOԌ��)I�'���\�_�+S����Z8��4���ʡ��	�z���v�_��Uh	���!�Pf��	-F�Y��n"���XV�M������PK�`�=��I��&�� �����7���ȁ�n�$b""�zל����Ӝ�72湫Xφ�?��b���;���
B{�dh�7��)����w�����%#��E5���w��<�#����Ӽ�oj�g���n�?P���Y9�dǼ�6,�Y��`Y��#�f��I.B+�/���l��ws��5�= ��}��$K�<=_�pl��!B�U���*���rs=��O�ꛞ'S�EE���CEQ�@�q��������I��Ȕn�3�|�_�˱~'\����Dgh��V�y�x"�#�П`kJC���E�����v�vT���/}��D�J����K%9̙*y`ض�z�RF||U��V�'���b�"o�`�}��L�V,l�n�}k�{�9q�Q�rެ��tp)`�e4*��?1�S&@�hژm���X�rK\TQ�;�a�86�Cn;�����i�8ǌ��٩?r�`[�L����2X�ZW�3��A����(e�Zu��g����2���\T  ����o��5�߫S�  ���_&Ѳ�?�Z^��9n1���A�����5@L��_p��nD\�q =+��)��͹��qy;ή���a�,Iy����1n���j����}(�Ӯ��2�Fe���n�ݼ���>�"ͪ0������s���Y�f��O��)�0�Ǫ�e3��"K�!���Ty��qp>�v�I�un3���_��q���͑��"���iP�{ǌK׍�������t{�r�`ܫ:C	�j!�>[;��_�����7{����Ja����wnζ����ݹ>��|��J9��S�0Q��)�Љ��x�vv.����W�H�`qd���Cu5�V�.����d��M�2}6��	�& "E�S����^ohu��%��X�J����d�6�K�h�[i<&��|\�4u�!Lbe�URWD'.sE���=O}S�W�#��'�{���r��x��G��B�����oｽs�n���a��DV��A�[O�������qq/\-W7Ma�T��&���r����_Q�	�hs��������j\�}��ɱCm� Y��J��.ehu�p)��ы� -�������N�ȑf�a�y�?�ܱ�Ξ{б��!��r�ڮ������/]�cu�1��)W����$҇nT����4գE��]�~�O d��}�g��{Q�^~��K���@���"i	�@zf��\�������b~�Z-~d�o�r��?,B���Z@ aϺf�P����n�	��o��<ݼJ0PW�!}d�M=�')�4X�r����6ozj��3���Jk��>��r�̓{�j2���ʍ�O�^�������.�7�Ԛ:rT��_��kG�<����؆��!XN
��s�7DK��z���:?������<��e\���6���'�ѥG�v���>k�-��mi������#$b^`F޹��ݾ`��eQh��N�]Ec|��v�ɻ�X�Ո���X�-(L�\��^�눤�`0X�-Lx/\;%�|v/�Y�wi�6�brg=�|=1wt�ȹ��}��Z��'oQ��p��5��X� ��S�|.��S67npi�9=�X������2�o�v5�k��f�
�u�	H�f�я[q~�%�1�|�x�}.|F,�{�]��'h֕(�6T��1��Q�H��ʚo��}��wF��S)ӛ�-�,�K~���Q	�V����58qa݉��^āĺ84��>��e'ǜ���7@�L'�ճeM�6�"~�Қ������c%G�����<�� SY;�3l��k��n��x�v�:�y��}������	#���8v��Aȁl�\^���k@C8O�W��iP�c8?ס��ͬ�����3�8�1�N�(,�����#@%�g�����_ƅ���@��W�� n�l"r)�wW���/ע{��!*�
̋)��5�F��f�ݢ�1��!V˷��V�r&��Fg/K��ӄ�����ʾ��n�J�Z|S�]ЇȆ�*��Vۄj���X�qؤ}\�/��%�4`2�}��l�h�����������'�ePD�V.�׿n)<�Ϻ饐٩Lw���b�r�~_@vϻ'��)M�+m���Y"���k���-L�q�O݋ɬ�"}r�ja�C����q2�(���r�}��[I|�ٺu���ka��_�|�^���sXwH^;/Q���I�Z��+�M����R����ʁ딻�`�c�5��cyA�Ϸ9{��-�6P/���M�	��|��{Q�Uec��Jyo~�f���r��z�W�T��tUgcx3� ��do�_���g�WQR�R;�Ď}��hK�t�7̑ٽ��j��j�K4��=��;��q8�,&�j=��c��v��5�⸭�U9N�m�P��XE��5�z���F7|Ŝc,�i!ox25��&]f����]܋p���j�	E{�h3*j��w˕#�2�g���u����v!����2��.�g�,q��E,/�4�<�ݙ�IjX�t����������l!���E�jyU���� ̮wlKq�Fs4��h�v���h�b����8�Z�E:�r���a��Q�zʲ�-3��f�Xocz����jr:(���_+s�c��!X��'k�z2e��f�fB��+��c��+��ˮ����/�ϩC�tě�af�cF��� [G�����dI!엯�k-�x���S��z�'��g-�Y��Ftb ��R�t�j��"�=b�e��ሢ�
��Y+���~^L�j�%g*Ūz VB@8�qۆ3�/�Xu�}Z�.����X�kXv��>���z��G�{l�ҁ7�q��g�ׅ=�6k�,&�\՝y�QXa���a�B�Muɽǲ��K�N��v�q�̘�����/*�*姤��KKr�2���- 
B�3��ݿ�kt�����/]���X�r7W],��Tmwb�Z�~�7��'x����c��R��\�E%�L[힅��T������>Rv�t�[1���5'{��?թ%�ic N�o�V�F���Bl���;��У������"С���}�\
��xMM4�%/��|��:��fKeqX��D_k��� 5����p)�1RD�3�_��A��j�պ`�_�5.=ZYY�xW=�p���~���n���E�sW�s�C�Z^���-?X�uv���|k'#����gn�8�7�MC-I{vi�]�iA��s%ļ��(ev~�Fނn�d������Qg�?!�ķ~s?���z��ֆ�P�9���S�?[��E�12��)U�]#�n}/�vCN���U�֗�
�;֭o/?�^o���3n�q�@r��,��5�0�ʭU	�
�`����%�rn��x�b���uE�Ȭ|%V���}�p���O���a�z�j�W����m�
�g��e�%����Ke3��5��yĚ��Aq��؃/%�-�_o�^cg�g`}m���0շ��>6�R!����2�K(���ĭ�*P����`pZѐ2���������j%��(�47Ìhz��!����I�gw���V�k��(H=p�q���?�KXv�:�a}�=�T|��>4R�9as��&A+���{�݆�^��aj�U����*j�xWN|/���B^*��� u.T�q,��<������@J�p�T;Ȗ�����=vZ%|�_d�t<lZ+y4#���7����SO�
^s?3.g�jRs'Z�C��B#�����^4	Q?�=5Qn�;�UP��q:�+Ui˔[�g�W"��̘?��<Ş��Z�i���|���2��r9ǜ��Ŕlz8������6*��L�1��bA�В���5q��ֆ��݇FL�~��L�`���_�1�F?��7?����'~]˖a�7��7�b�0����c�>�;�J��i�Gf���-�t��q�ϭ�Ľp�~��}�n/$N?�V�;׷��, j�C9��UO���=f��,ٮ��i�����¹�Ae���T�G-GН�L���Re�(HK��2��X]}�p�wf�-Z� ���N�T߄��#/���/�g�eK�˫��71i�ƣ,�"�� s���#��=7�/���[�j��BO����f�+ӳ�k��*n/x9������떺����uDTdF�����F��ә1WU>O3���	k�_oh��/CZ�z�%����Tţ���_�E��n�t�� ޜ�P���"�!3hb��"C�w�����sF�1@�K�W�L��kݽq�N/�b ����/�C��s���nCi��_��δ`W׎�&Ep�p��k걹3���۲�z�>�R�����i��g:d)U+�i�a�.v��H#��l�'Z���B�+����pf��&�/]���z��O .��
Ep�c��$"J���b����P�֣J���}��w}��(�M��`��{pa�Ũ 5k����9�n H$�kL,ɸ'�����S�����aViN�w��*��@��SxWz���^3���4,08:�踌������꥘��H��������!�a8
��ouK�e>�(X�:�w��=��V��= G�K����'}od��6m��8�;�b�E�� �-�4f�̜t�|Y�4KQ�cG��v��6r�Rv�Ӡ�ԮQ=� o3�й�@�@*$���߂(<aN �_��Ш�#?���w��|cj�w��M/��H��j�G�j��0��~��!8�����4n'[U,��^�R�%h�PwYK^>�`(�������T:M~�n���;��b�`��8�h��*�=�ꀾ�f��Er"���X�x��6���3B�/�%��~<�)�a$\��/���M�;�a�֗�ɣd��Z�m�5����8�\��SK<��	ELT����=dk�T�u�̣E~��% ��(
�%���py*��Vj��h��r�G�r�Vb=��qo�k�ޑ��s'r�����gy_Ќj��[������9�-��D˷CZݍ͈��Ħ��o��ͦ�操�b�����ćb� 8��I_A�F�� � Q�O�l�r`7s��i�ڳژ�,U�7�Y�_�r��d��<�:v�P�.���l�Z�O\� ��9h�Fm�异���V&Krm���ȷ�Y�! b����47�K1l4h�2�3�Ȟ��.^�V5+ˀ*�k�� x�eb��D�<ܰS�;f����ݫuЕ��~��ӗ2�k�5}ƊR��f�~�����`���h��|�H�'��!9A���X�x"�5�	���`U�c<�xԷ�V^v:��栬�L����-NX/n��#�UϬ�bu�d���@���ݎ�[qep&�Ku�S)üb�����P5<���L���as��M������'���U��3ŏG2��7AW("����ٯK��ag�b�u�|�X�A����nb"gg�1u�!�DIݑ4%�!��f���Q��T��Wv(��d����N��b��U{�X�L���G��{��'��!���&���QMt�h+j��f�٪/����QXK�=�Ė���Ȉ���U�3�<m��⿗�+����M�WU!ۍ[�
�ys%j���o�%3�X�����o���~%��h?SX[!�(�s�Ķȣ�F�m���-�*�޻�+r ʀ�T���cΜ���D�R'|C/q
��t2p�v�<��6� �����J�v��f���;#15��.�Ӑw�Z��(��I^D���r���N���Ҥ����=��C�����Ư�%c��1����C�r�cS�(��D˭�_�
�\�G���v�h%������ �/��7
@�7x�S�@ׅg�}z�?��Q��D��]z�Ђ������!���?{r�,s�^��1E����7@]�o:.�Qn&cY���Dr{�Ù.\jIU���/EX��y�|����3�+�/�Gf�,����nڵ,��qf �ׂKu�*��{o3�����O��{O�����zq��\.V�?����k��ꬪF�{j�.`?f�*M%^��u[p�4�U������	���a�LJ�m�B��;X�9ǰjC/�*P'A���S��X=]w���~|X\��a5�o���BӸ��7�e�nUN��LY_B��_J^���j��S�F�g�錃A��k��*g�d�SS�g�,*���?�����>-�����AZX��D����%G�O!Lɛ�A�Ѷn�z�����*XI�V�E���;���T��K�V�%!P�e�g\��s�/�����GV��+����Ԕ�\?D�$�B��nn���'/��U���ȩs�����V(�?�����H��
بӱ6�P���Y�6���#7���bP�{K�ҏ��6�i�Bm� 
�Vo)ON�7��� ��� ���(�L)H�U/�^��Q
AO�iW�Y�'K01I�&��O��^��3��;���G���Ws\�Q����40�0�-;7]\��!ʹ��5j���;���vZY"��.o��9/j��NEE6j�����OM��Ÿ��Q���t�N�A��Sa�0�z�c׊Y2?N��8�x	����?V�31:r'G���	��3l�� "��F�D��&>r��W����Q��mT��W�G2��§v',튚�nKڽ)n_ pR�m�gc��n5hw�T��xiR1'�B����r�<�ov��MOl���~CϚ�<A���H�����5�g��3���f�q5_#�F�Uj�p�{VIB��8��"p{?!9�+���f���v�>`�s��R�@�[N����3d���/jӖ���I/��fs^^e㒁8_����<Մ�6� 8�HH����_v�!�*DP�/�|�r~L\}|����2գ�+�ჩ�9��TV^�f`�q���l'R��?[j<:�ʄ�
G��î��0��jS>\����O��T5붕��gC���oӟQ"1�n9���"�VX��ɇ�0x�`��4y5���������ˢ�k^� [��l��~�/p�S���-+���7\�|?r�V-��;9��[Y	�{7"�1�ׅZ;wy��!�KK�{p:������(���ؾA%��iI���¹�M���|�p�E�ؑE��3�K�U^AL�c���b��1G��_f�Gh�a�ߜ��'L/����FT-O�o����4:�"f,�v5�eL_�w�9X�Z'�y�Xz�nk�86��w��N�-?�g$&`̃��U�WcOJA�kR��7d�'X�Y�at����:�Ծkp���bc)w��v�e�S�PC�Nm�*atdf�N4�k�m; ��<H��@�����/j�0 �_�U��LW<� al+<��b�q~f�bmNL[��)<��[V�޿����m��}�J�\Ȗ��)���nY���`q����֙d������pnAǔu|��@k�8���W
S��7y
l�F�qE��F�sA6)9]���6�F���W��K;,�U :ǖ]�{��+�?�+�HG,��W�����ۥ?ױ<n��i�
��[ݵ�gJ�����Ѳ�0l��R����n�?����Tޣ���K�PU�5ʚH��l܅�k�\�mTyRՈ���@�J�fml9����Ed.� ����Q���uX4������魣 �mnU���w��Vn��~�c.=�:�-[�ܐ`br�{	C���Е�=�K��@��*��mT��j��y>M2�J��I�s\/>R�����]-k 6|--�&`_��u�U�5��ʽE�S�ק��m�ODn����R� 򾧫[�Kq;�i[+��R���~�&�]�zؓvC֙��!h�>�\!L�Ղ��w5+R��t�O�C���m��s�����'�W���ʭ�8��s'kpӈI=��A�+��o� ��AN�[�As�Yؕ0ְj���D����i����?�Ҏ��I�7]�1s�P�e��4�����b�˵qԇA �+��������Y�q)d2�It�{[X�9���c5%������1"�=q�݊�{���*��K��W8���:y�y�.�x�H�����{;��>1ͨ��0�9�W����E<Qp����{IK�jJZ�Ӓǯ�-��=z��):j�}M捜ͥc����IE +}0�J\uPҒ��u;}�D '���3��G'���k��3��>�e��,��䱡�9r���(��(Hi@0�*���, �ѱ/t��=�iN���ɅY�f�𷑤�w����ӍY�zB?Os��nM�%���'!�L��	��lJ���耰�O�d�m�qy���t�'	A���آ����	�z2���e�l����d��֏��^+�{#)���7����:�L֧�۠JzÏj���i��q�L�R�q'njDD�ce�z��ԏ�{j��*ukwK �g�S܍4����V��c9�[�X�I�(99 s��������ӳ˥0�K�?�����/,�_� �g��вi�M8^�-7~������KHI�ȝn�v�P^i::�9���Pә![�_h,��B��7��زU�9���vsK�f�=)T0��zl/ݤʪ�R[`�����h���b�&�p593<I�>#�n�bC=^��B5��3��`�����R����L�}C��4��� M��_�_�{c����2\:w(=L� :�ĔQ������ی�7Ъ�/PU�1�����] ���,�U%bF��Zl���㳲�x<��� ��|�����ڋ:Ú�_���"tk6/'R���PU)_��g��8%eOY�����������ˣ�+��������?|z���'�F2��H0 ٕ�S��øv�D�5��HH�;�xrȧ�	�K ƞ�L����[hM\2BQyT�Y�c�3��6�H'v;*�g�	f�"�3&�	�mtٿDN�.��~u�qpf����;cƶОS.p�E���K�=��8~�;��n9������`��ɦ�u��:u�7c���{son3ވGJ0}�0uz�����KGOi�Mj����4s�K'�2��oʩ�Lb���4)'��"a�L�K*m�*'�tE^�-�]��_ߦ����jJ��c�����}�^� �Q��NEA@����* --6�G
H#0F�4��5���������9��}]��;��r65u�t���W�@84��`�,�`!j�������u ����ɪF���O��&X�Z�{��r�3�8�_�6��R�nY�0ft|����6{E7��� Hn�9��:r���˒�ht�����A�( gS������1�;���������#.��O�؅!)IH�y��:�2׈Yg�]�
l�8ÿ��B�K�jZ~��)�GT�ӡ܂%+R6��9�Ivܓ-���S�����>�f��]��#�>������$a��MiN$�k?��(�e.4U��9�ǝ+�]��ҹ��6'�r���[w��2/bAp��f��|�����x��A�@��5��x!���Уd�dT����� U��A�E�$c�^��-ω*_���p���f�b;d4���θ����t��\��?�½���`(�A9R�oK\�	��%��Tx<�4��\��Y����}�Xc�6����!��W��:���g_®�"���<N-z:E�{�0o�q����d��l�y���rVSܩ���BWח�	�{��ǯKfe�0�7�o�*�o�����R�V�]L�6<s�ˀ�ΰ��"���(�@q��_�r5\��}6�Uk�Q�?�f� �a<>��i_�@�@�<��[��m���,L�Ll�A~���O����\#��W�o���J�cm�˾��?_d�a�+�oQ���Qb�{��%!xx�e�;������f�pm/e_�_y�U5�gD�"^�\�堉̨���=���RD-�8�R��m��>ŕB��9:��"Yv��%ڼI׋��ع��:����|�(X�a:��sVJò��s�t��"���8�s�LSV���f& #�:�L��-�ʏ"Q�PRV�A�/���� �/0)�u�X�u��%�rce�ga�8nPG��:��y&��� #�<&r��&�f�{�b"9�4��	��ߒI@�ʚ�j�:'L�]�a7�	��}ԟ��RT?�㯍��T�&�rԢh�������zsmO6"=0�J"���"��ASz:6K�v�І�oܓ��;7K�R/ђ��Db�������>�}[�C��wPz/����ݒ����ۋ,�Z�W�r� �	h���Z_��.�l���Q�K~q26%�k�c��z5���ҲGu�M���;�fi�4._��l���
�Xl�A`��8� ��c�/:�(!�OF��*���ǘ|�H��$_R+�	��n4���*$d�w��ϛ����F�}��2��$����!�a;5۽�R������>r�n�Q$����������S=v��[��Re".c�B�JR9�h��F#��I_������ʩ�7~���ҋ��`���(URVN�[��ܺ�Q��TJ���Mn���i�40����9�Qr{ͩ�Umڝ��qL.r����Ԇ���w������X~�2��AkBl���>!]6*�<]D@*39�X�k�!q�!�8��2�������b�b��fjm<�V_/��/�)�S�Ȥ���Gz@���T�ޟ)�\UzU��p���_�`���Jc�s��5��MbFM���RZT�$���n|I����&k�N�̦�x����:HMzњ��g������B����㺵��*L}��Ě-��+7
�ءӥ�]-k<7
����JC#u�eҭՌ"S�e�<�����K���Ͷf�="��l~�Ĵ�ӳ�?9hSI��uY_a��QC��c�1l�8%�Ùђ��mC�Ò_�^�f���%JaU���|kyZV��>P�K'y�-~
���B����¬i@���|�s���\UBK*�0�F�}��������u0,Z�*Q���N^���1��N�.ZkR[�u���L_��_�_Wt��5}tƐ�[���C1]yT�HŨ�r���u͍�0��]�k��:��c
m�������%�x��=�IU�8N�B:|�@S�x��wF V-��%w��#�p����3�^���y�WT$��#��06݉o�Ei"O��*�R�3�9|��j��lo��[p�����ʟ9o���]V�&k%�^�HY?5��&���ؠxt6O�?-��:�S��Ǵ�8@���W*l ��w�5�IKd�-�q�(��-p��jw�vI2`�َK>�D�!A�II��;b�7���_j
�UZ�a���7����)��4ɭm�Vٗ٩��y6�7l�(谞�§B|��Q�Y!S�H7*O��:8$�!��7�ڟ���U����D�o���}�,ub-�k�'�oh��:��8�І z4����<���j�q�Ya�ٯ��%|hD��c��鯎+wӬ�P��T�D'
zC�K���~�m�Ճi�����X��빜
���SCi�� `�@�i

0�o�åڮ�V�I�ORLO%[��Zhk�)�l&�:|�yRº8Mݖ�(IF���}V���e�M��'�����Q�`.e��z�r��W���JyNg�kE�7x-�h	���G����}�X,�=:{T3X�)=5�}��'oӘ�X�&n;o�E�7(�J��x'�[�� ?�������D0r�?������F��|E��EC��];¥~��>Ɏg�pz�`U �׮�s�z"gm;�6���C���U�$�5��{<.��r���|y��(V�z��_�	{������fvX���A �[�$]9����y�
�J�g����?�>�=���^��W�&U���?cA���e����M��7u��.���U޵�j��kT62���]�el�nNl�MMK��^OD>^2����<��uz7(@�Җ�$�E��[\�`4��sƩI{{.ߞ�	+�,=j�p?���<o����|X�}���?���@\��􎷣ZD�o��7�"mi�Yd\��R��G�A�����v\���gUnv�և��t#��i DC��61e�<F]��8O�S�>z�s.e]�|�[O�p�͝�<�ӂ��$]$鑈�J-�����3eBȞ��<ChA&�-�3��9�_��1�Sc	_D�i�jW-;!a\�R�!\��6�r��6�R��u�^J����'>e$u��k�>RP[T�j�R'X�-���K����a�����}��"	�������e��uD��,ye�������F��V�m�Y�8ឤ������6�փX��i��b��f��iW��T�fr���N����P���# �������8ں3.^Ќf��N��K��I��2�vV�--i5�z*G��K��nO��JJfS�TZ��i�F-&	j�����Y�"�ѫ�t9�;�(�b�>��@n������b�%�~7�����s ������k�"��a�Kz��V�l�_�p,��w�V6&�� ԓ�M+�t�yvD��H����*��$3���z�/VP��4��M5*�!X��n�12��7���j!ۯhz��*�v�\�������g���
��e'yPv��3��q����Us��;1?��k����W��>@e���:y��а����5��/\9�f�A�jɏ:���OU����N7KL2������E,�QX<Qw]݇��/������4'�G��eO�S<򢞤�4xIVi��Gv�_T�N�/��<�p�3�GI����j7�NN�U�ND���t��yq��צĪ���ZC��9Y�ւCS��"�[����?�iR�A�5����Ü�:���L��c�C����gl���|�.��ζ81�)P�yu��T9(>߬�����1����7$�N�s����?����s���=��|������g��N5�" �I�7��	�7���8oZ�g�j�ǝ�&�R�T�l�i܍�w�g����!�y�n6�u�$Į�9�I
{��{y�#��h�5��#�U�Q�L���?��*�����uw�����`*����yW���T��5m<Q�����/��a���ݵj����w<J#w��hev`�r�D�� a�|���>� ��r��aT�|����.΂�췩��e�5
���!���:��b�쳝"P�v����T��aU���"���Z�+Dk	7���_�I�8�D����3ix�%����V+�!���σ|�C����K�:^�;j `�:���a�7�w�B���.��>yD�60N���F�?��w���5J'�������jS�̃5َO�3���]߿2���ǖ�+l�Q�s�;��:@>��h�B�}V�\������k�SK�ӧ���n�ɦ+o��W�Ig����]�\U�7����b�>m0?l����7�U�L���&�����9��`mk±�w��'2^�i��n��d�����Nw6����6�E(�-B��$�})��
���]�n���}'���o�>>��E�-�(�p/=D������¿��ƕ��
����+I`�AS����zvKa�/0-���~\�\1��xߢ��'�T!���29_����NJ�ޮ�f�Oڧ�=��H�Z����)���O��=
�F�1�$�d�X5ͷ�o-h�����8�1���}�.����KC���~3:���:賂��%�z���3����2.P_�ܡ �e�؛�1^K�K��Z����c"�C�E[uY�	ț@'F`!EE`6�vRU�����N:�u�����ƙ������1Š_��|u��H�QMM�T�z�k�L�W���J��6C����Ǳ�2I��d�,"����~���g�T��#N�`����?�Wԇ�`���	O�����ģ溛�ϑ��Z�}2��g��~��m�&e2���;;v�%=S7�+ۺf���5�F��-���	L��l�v�ëm2�&���a�r4ɶ�������n_b:��H�y1�BH�L\�����L��#>��1_+M����[�>��x�����V�^��];⧨�J�'f��2�=1
3�\��d�U�σH�K� tя�`::�}�K��榈+^l]1o�2�-��G���g_`���4��Q����x�����b��}T��!W�yò*r��[�u��&�2åoa�{9ԋ1 C���pST�M���س��+*������q�.�wĽ�[���Vc�?��|)�5֗Q&l�_��H,���☪TdW���鳲�����0��>����5�$|jr�ͼ��Ds��)���G~��f����җi|�����|8�$6?l�A�┛E��Qs�� ���0%1G��s��D��>QT�O�#�y\�N���v�"�ꓚ�O&zCL����w��j�a����ԯV4��U��D�u
 ��u�)�x,�7�n�X׭d��3M����6�����BY�}�\��qu3��&�("Թ��3��L�0m��V�!��T��x��8�?�]�a�oV>�u�+$f�̗���89�(O`�¹���ײ�riD���󇫤��>����@#e��z(��L��q���g�B���e|+����QQw!���C��~[_�=��:8���KqEq����'uc�Z���..��c�$6�M��ٽhބ��.�@�j�y���s�A=�@�g�
�>Q�@�:��'U�)q��:c0�L����mTv��;%��5�ݎ��-�k,�YKIY�^�eJ|E�9W4
&b���I+�;xӶ��.�w�x�m�/��5t��H���aI��P�y�HPA�wV]��+͡<,$�!�k�n���8���"��q����4�dwm'���c�T�W�~&a9�KۚU�tVE�J�=�y:���1r�%����f�XėI�'�#��w�P������~��_�Wˬ��$Ɖ�9���|�Y����T�|�V�B�H��jL�I�:���2FKTfK���g�@w2������=��F^�L~I��C��l�K�����#�B>�C�h5A�-RTa]��3�����ⲣve
��98�v�U42�韗D}��%o�x(���+���.�ĕ+�}V�F��I��7}H0�	D�mf^u�7�$jC^�J�|dk����,L>l
�\i[�����]0.|ӁY�I)u)�&�C�7*6kf��K ���s�9�m�s�͢��}��K�<_��$��*� �`��7�nkoW��濼Z�_���oӓ�jDUX�����* _(K�l߸V�n!��9���z>8�O�ͨsw�N]��U�Cm�C�����A3�]��x� I�_4gF���ݙ���*\��ی[Ww�A��	��ˡ��9_�KD�����&�}Fu�1�_/a��Ru|l,%��%������_�=�n�c�{w�6`{�7�7,�n�n�k�&Jg��V���ZM���O9#�0��M�ʿ�Ĵ���� R���T�����)?�ؙ-P��g�3�� ?��o�ݥ�G!���ϰ�3	��O����۟ʋ��&М���wb�&����+��V�D�$Z賳��]n��SdX��Μ�
�GѬ�[���S�F��1�J;�"���3p��ﮐff[��͍��#n~�M�k�̈́��)�3�m���He��R�ؿv�	+�Wz�a�]��o��ƶ�����5Mh�`�h��x�3Q@�$�,��[���;�:�K�<��#4�����%uѫ�t��4���B}�܋�a�+�\!`�C.�݉�ڕ�,��N��x�-W�-���o:ˀ�"�jZV|��2)����X��Q�������'X�'�A�t.���b�K`3��o<�lnM/Q�Z�͎o�+�$�h�S�7�5K�(.��!���X��q0	��|!��2Ð�l����:Y�J����>~+���ٝ��}q���!���� /3o�pR�m��k8߻$>_ej� �Xl�]2{I7� �\��9���CPJ���=)�v3�	��ԉ�~�:���@�h3�Yȫ�>�^�_�I 䙃U���z2�T�����H�1d (��8Og�11�M�����[��7 _�FF����p7�רQ���p3����Eyԍ�4eM�����^I�/���m�Q�N�Ö��t�s�]T���C�;������4ű�\Kpx�O�Wʢ���a���dQ8BG�#�~Q�9��E��Cթ鲱ޜ�O���U���vl��L�A6�7d6�~��^�'�A$�ƝVY^81&m8x�N��\{&B���>����7G����5��v[���*�M���qㆅ~ܯ <����TC��z��4�^;$��q��iԎO[���?ɬL���0[�
&��/�G�vv����z��a�y�S�DeG��DW���)�����9K�x�t��T��UX��l��
�A{/�յ���t$�"������>=���?�{
��o�υ&���..���x��3�m��i�(����ꜜa���2�}�dR+���(Ĉ�SR��,��K���*E,%�S�ɫ`��nfN0�;y��l_���
��S�7�;RB��Q��BZ����ڂ�DQ2a��^���Jr-�;V���c�ݖ~��E~<���PL/��(��=��k�T�<>ؐ�����(^m����b)��D��TN�M%��g����`{$-MR�ݻ�GC#ȃJ�Y:`��!�D}Q�\�;؈^;l�mR��[s����:�mu�C�ۺ�e-GGX	�F�����2*��#��d�~= ��Hxm��N���!���	Ĺ�9�V��V2frziGWzl�D���=�I�����:뽕ʵ6w(*LYw�ag���<������ņ�t��rרּ����ݱ�C���`
*Bۀda�?D�;׉\μV�A�PJ��'%Sd\i7vo����	kDS���X������x��3��qƖ��ǣ^H�(�e����ӟ�����W~7X�?�5<��gj��޴��M��3�4��]�T�Za��r���P��f�x_x��9_�Xh8���\�ϴľ�~����_��K�	a�|l�_\^x������e���V�	����俕�Ư�S�)5��9<9[w�o��m��B�v����S��{9�|�?���}��H��m�+��W.�֞R�r�&�z> `'�u�p&2P��&%���+i����@#'*7�#|]\J����%1y���UB�&�TI���s<�]ȡ�x�c/��m�����֍�@�ԣ�O��s���/27�����f�#R�e��=W�η�4��7e��M�a��/ۦ�Qz3�o����'��z��mMS��-�܃�wD��̓���+E�!�ƫ��t͜C��r��oNTu�khDrrHI�.���hd���8�rv��dA�?�����}�y�uǧ-�EY�[��8�l�����am^���G���+�(DxhD��O��,���ޤ��y����"��v-t��r��*�>�v�U�;��n�C�r?�m��7)I)ޗ��2�7䍱����(��wԟ�~N�y�U�#�͋����K����"kY��z�a��!2U8B�B����?B�^4}��ă�^Z,�<[��:W�'���H��YՌ؁�V��ߕ���v�Uvƺ��
2��PD�^L�}�jtqZ�T@
�����Z����ʨ�5b��}���~[�$܂-�Mtϫ��`^��Bx`�=9'��O�'e4a�9���"  ���Oq�vil����/]��|U_�Ѐ)��Ѩ���DQ��r�f���:��Ŝ�F���[7��ۘ�+Jy���m�_�f:�����N��1���/��'�R��v�v����`����A�oޟ�ڡ(�	R����q��zfB���¶�,��M_�G�)�V�/ㄽR�t3����s�iڦ���;g�����҄�M��p�7�����L��}�Yo�p �OH�q�M@*٤כDғg�¹���}��O[؈/�+�ׯ1A�G	r�"c1���m1��ʟ��R�J=^�+9��װ���}�fj09G'�QO����kd���`���tȣ	H��uD׸��D�;;5D�	I=�U+�uޥ�o�d�z���4y��/��d瑭#�q�j�Q}0�~`2$N�Y�Ii,�ֱ�dԹ���'��##�%}���d�[߃�'�Jis;�m�K��?2C���R�d?k���W�v�EZl�Ȋ$��=|�4��H��\�H~�\�;�FA*�C������\(}��$�6us3&&�b�S�o�<�3_e���$�#�����ա����L�(�I�$�s;�ո���_����ә���
����k��1D|�T%��bٸ��ިq������h�F�q²�Ҵ_
t0{F�rҬ���BK��#���,��Ù��!^@e��j���l�FW������*��g���=���:�sY@���S�)~Ŏؽ|K��4����[B�W�CZ+�����K�����/�6�/��T�����c�s UWuP�^��B �����M��T8Dt�P� �H��&��\��us��RZ�2l�L��Iy�[�~����DЀ0*���G+>�L3rv���H�8l'�����=�Ө�(���L�Hظ� !�V��3o�)���X������-.RUx�E���杞�e��S��"3;�����0�B{�"t���|qy�[�}Ǥ��:�S}�N�Nw���!*JV ��ڍ$rXO�|�w*�d9������ǃ�>�댿m���[	��.L�\tx��aO4���b�Ґ�'���1�<���ࣼL�:����orI����DK�9H�1�Lί������k��Y����ua�M�������8��v��i�BB��;B�%ލ�b+ˣ�o�r�}�e>0∎��5u�)��g�+YoG����1N���:fB��!�{0	r�〢�;|#�|#[W��(�ܽH��6��@��). ����&&��K�����+�z����'��yQj��@�GRۢ;Y��-yXE����B�j��D�Xk^8m���I,5P�Ra����0��g��m�͏V2�>u�ʣ+�/��f��}[�3�L;�"Y�6���U����
j�Hy���p�d�&qV-&j^u[�ie�v���iD �ʴd�v;���'�0�&l�:W��\b�G��D�j�H�kX�E�l�f�V�2Sݲބ��l���v��GA/gh6ꢫ�3���e��â���آ��-����G�'�ag����)߸�g���5�ˏw&N�wI�>#?[舚�A��3D�/�­?x`��Ӗ�:1p!�g�j��ک���r%/3f�Ԍ��z�_F�d���@��$����E�X9x6���%&4s�`ֵ���:�L��.9Y�a<�N)x/�*l��Ku�����>����ŭMb����{l%�]� I�ܿ*9Ձ�&��_�t�IL2�5��#��e��yQC�Z���fG����䮼����2���Í���B�~���? ����A��%6%�QS ��c�|��2�K5��s:S��&�}RM:Rz|�zt��.Y��]�,�mv�Gei�'V�;kh����x�Kx.�\�Q��<&k��ɫ3���Y*��n�U�x�`i�K�zl5�}���ڭm����s������v�gl�sŶ�i�V��������B)��Z�PEw7�h�s��?�5�����kq�8���b�ʁ�w�Pw�"W�� �I�����i	�)�6^�k��=��u�Z���I�A����0U&&=�q�B��E�C�,佽K�Ͳ�(�14Bc�-F��G[<'��~�.�N�rre�>g^��KG�� �Cb[�;�P6_�z��A.��۴�х�deƇI�"�2Bʏ�{��e�L�魷b�տ�B�J���z�8c}ٳv���3Ӷv�u�q¶�@�|��֝�����e�IJ�Ju R���E��n��C�m�צ�������ȕ�VD�t�&c���.���g��z�"�S��Ls��ΕUt( "��u��7�ѐP�p (.� �J�UJK:!�o �~�1��_=3���=0��X���qNHB.k�G
J��=�Pc� $0����|3ǽ-.�먜&�T�FU� 1��zii
P���5Y���I��S$ʰ2��`�U�o�� üH���;�@R{��_ȴP�iv�L5+��F���sY{�93�L�������V#��ή�E��l�Oh ��N���Q�t<k��W�ܣ�h
��ARD���G��������qʶ��[���\ӂ�o`�~��|�����PG,vm�G�Z�t�k�2�lK|y2�7��ɝ���Շ�����?����:dgq�W52�pJ�q
Kg������+�����\>�`�����s��&����"�c�,S�G���?�H{�۟u�i�5jj~��;�M�w�t,���6pL�ߨ��94�O�|��}��)jW9yp��G|���kv���}�8c�>�F��7ũ�(�Cqm{���7r+@%�&�G<?�&�*]�"/O�> j���Q�޴�@8�/��Q�6���x�0LMI�N1��3<w��I�@��5^��i��вno7�M���s�{����	>��t_#م��Ks���.6��M}�*2�K���i��%ғ�	w�=��,�(�Z�ܵ_�H�k95~�� ,2��9����^J��b�3.�Rr��P�OmO�:$F�G�T�'�x,j|򥡫�h�p Y�	<(+��0b���+�B��BPU�.b ���`��fX�.�@C����+����}u��2R��)�M<?��CP��m����H��ba�jЄ�7��+��U@���L��Y�����4�>=)
�۝{���È�� ��J s*+G���0�z��ǲt�EOYۄ|5�,�9��'����,X
��\���=C���˽)�Rԣ��"����(63�Jk��V�s_�����V��{����ks]��2���v)��]}��FH&�:!Ȁ].��s҅�yp�1S�ֺO�BQ|����%j��Mȧt̸OOd������e{���8�3aǁ|���d̪�GH)�T=���I�K&y��j����2���E�x���~�QĮ�|��1Mo�jՌ�����&�[�u_��G���l�!�w�0 �h�c��j��_���ؗ9LF� bp#C�M.�ъ��|��U��N��i?�05�� D@���(N�I��ȉ��o�\OW�^ե��2�6���)$�LoJo�����-uD4��+�l�+���!�#��'pFӴV��e�1etӤ�I�������RMj�t�/��$*!���>4Ea%�[k#z�#�n��o)�X���
�@�n�;R_�ḻJ�3^&u�Þ���������z��)�h�"��}B����ep�2���~��\���"��`�������m�s[�)qJ�@3w�6�C����#�ϽZ�+�},�U�ֽ����**���k.���G�ۓ�lc#��93��+/ݍ�Q}��!��.�skQ!D��V�)9Q�Q&����8OL��c�2���b�~|�:<��Y-..�� s*@![O��+�*�����D��"S�}�^v�eQ��P��PW��C���I��j^ȭk���9�+�ۚk;ĳ����+m�������������>!�|F��O*0�g)P���+����}' I> �C��z΍���w�߷B�:�-,�9������m��y�F6~K$��q���ٽ�S^*�Y6^��~>h���^Y�to��I��ndG����\�V���q�*Sg�����ׯ>��(r����}x\ϳd"�Y;v1�=���l��9[ԋ;�S|ο�r���IJ�7S������G���06��[	����x���BS䀺ӜrU� p(e���ґS��A��D���/�2_>Pؔ�*�h��`�� S�l��C�A&,�܊�
���6�h9����w
*9�L�tz���D��4�r�I�Q��K��2���f��R��,I`�D�UVY}��|`��N�7��V֎?�`\�zdT�CWl�=ބ|��/Lk3���s<��O`Y�|������J�<[_�D�+��w��"�>��N�ℚ��v���T�{��P��5!�>v��S,�4�w�݋ 1х�&"�#��Wۗ���]Xd���L���C�9�Ӑ����]������A����,4*f)(���l^^P{��h�`j�A�̦��w����
n�5���D'�Sgw�ؑE���%���;@8n�`rf�z�ܬL�;�Ɲsք�$X�W�+�H>�xp:��9�]����}���%�%4mB����Gn:��/!S��FNjA�תz�$N^)`N�Y4���<Ӛ:]B�'��a��AJ4+J:P�[�s/^�?H0y��lB�v��?��vP�T��� ��/+qii�w�VTTP��~�������1D��k�׺�Fְ10�v�>\��Rl�ISg�X���p~r�-`����QT��Q��R����7-�$|���^�h
�q�}�[�[@m0O�^�-��T�F���C&x���Ip�j�L_Z���k���A�q}�x� �?�����{���-4ҽ�����-E��ĕ)����m�<��Guz\'�9	�+�u��J`�SYG��;��S��v�ҿ��oR5���2�TMk��:����S�8�&�+n�09N�O'�����4�kƯ��$ӛB2�5Vr#�1��<�(��Vt�|BYM��&��\ƶ+ޥ��Vu��H��Q�!aj(s�E���Ǚ
|'˙� o@HH�Q��s"m/�aX\��"��y_�Ae����w�(t��;��]IAȇQ4I�l��	���|p3ӯ�����q�3��B�s��Q!|T"��ZC��w)7.}��&���I}y����V�����D}�?����k~�.eϹ��Y���9f�7D��OCnR[V^BD"P�ޓ��|��D��^���h�?s(N(I���&��H6�q�{�|�n{S�ZP`�?�
��%�1� >߆Jy�"c�K�tO$/R�_�g6�u�V�c[>��4�i؆�7<�qsu��?�PXÏ�yō��㻖���=�ma�A~�=��=�1����b�%m����xU�ϵ�f��%��^S.��Ɍ���0憈7�5�g�a"1z5��dqm�kw[-��jkk����[1�x��3lG�m�wH��(91���S�C��Ƚ`$�Y�T������/��i��T��-M��%�bb��	C�� ��f�7�7 v�㺆��H�*鰎����)u�����e��D���*�`�����37��Q6��Z������rﲖ"����1(��v�c��*n��?��
!���`�W@�����3�q,t5��m@��8N�����nn���P���	0�=q␯S쇿���Q����rZ/Xds���(DT�:G�8�����S�Ȉ�ټ�7ēm�S�|�y���7u��i-y�1N��7��͌�BH�>��mj`.R�-x�ˬ�=���f�ws�q�����U���T���W���(� �abj��dr��1Q��V¢Ϯ@��E�UA"�b|�B;*EǱ�U�H ��@�"����ʺ7�M	{q������*%�8	������I�m`5 8��~���ؽ�RW���[���e�:���qG8h��G�eQI���Ô���_dֵ��e�*�g�~�����b�+V2�R��=.���©!����̐:��m{N�.4�Rxg�z�'��t�J���8�z̢�m:�H��8�L���t2�ǼEhro�0� u3�k�Mr�K �ux^^���B|��J��|�4�?-�D��c/���t+�6�)VZ�񯚞1{7y��?�{Lс��̿��RN�A�6�?͚�F�e����a�T���e$�8��l	1��a���՘�de��i����r����ͦ����t&�Ef��<���Q(��5a1~�[3�Ȇ���e[k���wU 2�����d���:��יD����.��[I�7>���h�`|�8�#$����V���F��櫘Y�hu/D0Շ�#��%��oQ��A�}�{������i��8�ؔ��2V2b����v<�}�>+X�;
�#�Q��mq�-�<���D�7o}9�F2Z�L�NGp���v��XT07T4�Y>��P�n'�}�����%C--�����"�[���k��i�TUF�ޭ9g��>����!��ac�V�w�Re�4! ��n���7����Z@�pU��>�t���B��QZ:x	<_�ŗ�u�E�b�O�U~
88�S2.��a5���l�����#���%�31�M���Vx��J9�S��:�ȍ�����X@j8M�1~3���Q��;�j��s+�;���qpШ�*��ɮ�F�3g=^�Q~�]`.�~���H/�`��K?��}Ӱv�6������z7V&3��������y���dL��}Ϩ.�K�d���r�����.
ӞV1+���T3x�<I謓�ҎPz�,�V�枷�v�^��ڇ"���/{������V�����{�f̞~����ov��vI��u4ؙ1gU��U5��;�:cd��+Zx�۟Vd�\s9Z��ސܤ���g�X{������dR@O���^#ϯ�H��x]�?��mq9�3c ���'={J�9cVoo�c�q�n;m�����(�:�����y³�E2����#MҾ�Gsl�,0�V[��޻�	�Jo�W�����ag�K�D��~w����ˍx}�nվl�:��l��J*2�/f�p���'w�}T�E�TU(�����oҊ��$�]�x�������l��Hο�u�}0��F5v�K��^Q��)�	0�M�-���U{�܇��6�/Sqj���F-U�uY���ۮJ@���ߋϏo���2f�������k~G�����P�iB�'��J�և����y�M�����ڦr�����l�-MR7+�	��|�4��qT!�Ѣ��Fa����·&�J,�P.o'��i���a�Z%&���v�_�"-;/5|� jS}�j&��;��}S�u��*"��3t�.��|hY@�6#slpx�Lܖ��b�H:�k�} 8��q�ׂG:�&�.�0�Fɤ��E�5���c��:U�d�iF/v8mz(�b�"�� ��Z��4��wK?a&W��"�O��6]�n� y��(1��(�Bك�>�,���I䆥Yj����q�?Rrc�_K�r\�?�H�y���ʹv^b�c�UZ�ީ�]�;ua����B�xn��X��l��p*����؎���u{s� ����؆�����~�����}�޽�*�{,�+2<�[a7�,W�}.�|���E�/������`\t���,��87'��t�8 �CH�͟<�V�v(
�RQ�C�D~CE��H�Z/@7��xy�\�0�ʊ_`u�F���6�I9��A�pI�~�~D�\���dRRT�7?�T fڳ���� xA�F5�cG��,z� �_r+��{N
`�^��y[]��O�zP���^��F$J=D���y��g�hQ��G#2��H2�_K8Q��8K�$:���I�ڶ�Q⊘EoZ��~Ct��	�����E��v�o�5�L�\(t���@i����@���h�Y���ӿg�.��g�%������y��0�X���a����X;�7׊8ˑ-)
�#�@8�ƈ�J�����[ ����9����%�����:��
wvwA鵵��s��p�Ӆ���qừ8���<NH���gf��d��Ɗ&��ʮ88MV�����1�
�Xd�k���8���G�h,@�z]:l~@������ڿh���t����C)��P�qT�d���P���o�:(�%��fBSY�!��R]?o��)d�>Ƴ��S��0 �"@�E���WC�W���Vf�NN�muw�a���+ �L�.�nk�&�P_j��P���2j��d2�о�h���6.$���ՓEL޶\g[i�QFω�b���q�]Nz%F�崦�D�M�_�(�o31n���T �낵��@5�,6��KP��T:���8-�Y�z�Cf�U��=�u<���3��̬
m\��J�Iʖ�@�s]W�L�sA�Aw=)ޟ�u�:W�X��!]O=�N����C��K��X�j������1��3��kg�a���=�������i����n������-- ����]� �"�������,],�33w\13�I�ho���?� �{g��k��&��W�j���?�c�j�������3�ǂ3��F��l�g��ﾲ>5��(�PS��]�U;wc�5cU5�L2w\�h�f[J�����=���'r��&vI��k��&/��a���g4^~���%�k��L/�o��'��ׯ�A��f�i�$*a���=��s,��kgA����)��?
b��ӯ���'sz	�<	����z+H�mˡ?��X0�=
�Mt}���H�=�?��A�����%���j,��w7���77U㥢�B�m�FN}��=OE U���,��#�MxLd�=lE&�03���PXe��qt�1�(J��~Ԟ���!�>-?����e6���E!u���0��+��֟$����s�P&!5fG쬏\���c������ǈ�c�O�\i5���8P߸AWS�ydFe�-Ih���#���Z>�pwo���U�����2���w
�X���h����;�5�?�f~�Jg��;~yL����?8�^4$��ܶ��lk�ު��My��[��T��|H�}Q�8�x���=n^&�^�]D�ڎ�oӛVqqq���w�u�I�%_�ۢ�P|�rH�p�#��͏"G��v�xkg|�P'7&����F��`pqo2!0��_����J)4na�<��xǬzP��L �FvKm����a�
�f�%OAA`b�kq��_4��
���e�k���-���a^�ߥAz{
��DބP5��
\7$pbLLx��z�g?C�'⑼]-K��Q微ѯ�Tv5�����[yT�eǕe8�p�]����4�O�pIBb����R�S?l�7"՜���&�q�D�J>VJK�<+��,"m^^URR���K��ۍ�^�E��:99��!b�O���#l./���Dt��@��bFm*ی�O�=����zq�(-��,���Nb�(�`�\��y�? S�;�S��w댊UYіdSV�CE$ĕ�౯�Q_�~�O���ч��>>>�K�������\Q� 8ݭ�)K>/�	37Z��,>*���< Y2������Ԍ�w`M.���<$�Y-l�������EQֶI,ħ�BB���j��>LŹd��-o `*�q�c�-�j&�c�Lͬ7�iq�7�(���or����.?��/�V !�$��1���G��E}P�Xnvk?����y����h5��r�͹����gT7��G�R=��}>G��#���8d.F����i��y�� ���W���+�a����{���rN��b���t����I�J^ЇGB*�j�,�~$3�lm��.�VD}�z�}tf��9��_���mT7��L�snL�3,;nk�=��[M�g�����X����Р������M�l�^�Q��vW3���4��_9bs���ⓘ�G0���Ec��>�Xjs0ڼ���4��x3@ �,��2J,��3�uU���X�usʥ�-�������}rk����!�������'�6~�����X{~ 5��$t(���>\"y����R/.�U%.>��k����}���4/%p��K�k)e|�߀Q_M����������`��s�q}z��S�l<�+?>Pp:���у���>`��H����ZF�����=�ے�חZ��9����tN}�?]�W}\^:Y;HR�4o�����='��������Ϸ�����u^�B�p�K���s0;�m��O��]��,Uq���w�Js��2�5x�t�^�$
]� �``t�g���ʪz?T\T�۷01)	�Pc����~�$�B�Bg��
�[J�W�$���YM�����_}��5ջa?����(�1�m�_�Z�5���쇹��m��.����Cu	W�Ⲁ�wr�:�⪪�����t�_QP����?z�{������T�Km�U�x����t��n����k8�:�ܴ�^���C41�˥��cE��F�J��9py[�x�&��� �2���)]��	ڭ$;9�x2_��_��ߏ�vF}����}I\:w�q�za��"wW����_h���gfV�h��c����0��#w����#}�9L � �vf��â���u����O������E���т:ř�i�_+pt�5�i��� ���S(-`c��n)թ9ϻ[c��O�JK�\;KKeF���d���{��H��qdx��!�|�'��c�W�_zK��Q}�z:o�v"�}���de}�Y�~a� =��B�e?2�%+})a|�V8���U�}�.���h������	 � -�6~7�}⃚��v4�w�����h�L(��.H(4R�2�GSl�T�u&�VXH#�ۮ.2�)��j=oY�����;>��d�H���IJ��򄃠��ԥ��b���Pްq����5��4:�#��sU��%x��O�qP���v�1� �����)��'(��^X��O�	v[����	z��k���t���4s��u��a���1!���n�� q͡ݤx'@+�m}�(Z�LZE�����Q���N�5���Z�v/,�?��o:�z�����@��0�C8i���.fx��M������f��d���5���皠ݭ��[#|J�nf��
93b��^�V�^�Yе#�OD��E���z��`��f�Yqa�~�������n�ʍk+:��#z+��J��?�Aˡ�v�+H�`��9[��J@�Y����e�� 5�)�-ʜf/����S6k� �y�K�uӅ(�M`-��U�w)�X|W��7�����\
�����'���Ø>Ѷ�^3i�'�_<�º��5^g1V�?�]��9���v��W�s�� �������}�Dd��$N�� �z�h�F�w����%��*HN �������Y'�O�ͣ��z��R�8��2
g��(p��/gp�!#K=�u�}�q`YO��j��R�����+~�7qD$������b^���
�ǝw�����gtڑ?��E��������kgf��eM���d��������oN�mTAZ+�l�{�iq�O�ol���=(1&�$�v�G%J���!�n�h"_^cJ1��O)%����J�!����y��}�*�5)5��#��}T~�n�֖,��%S�4RH�_;e�˅V؊[���~���������*L��Ƕ�	�ܘ .�c��fzͯU5Ct��������a���H�5�]� ��u!���e̀���L�@��};9���L��%�϶U#�qE�~aCpf��7�W�~�O��C�8ʆ�k�[�`:��cލ���9����]��)9Y�-X� j�������㖛�/7��ܷ�y]�鎗�o�g�rGx_�f&RyT2�P+�s�Vlӳ�̟m�5��y�]���{�	���(_��ڔy��Ge�e����������4t�m�]�s*���)���䂅�Ӳ�+�z�F$���z/j@t�����Yo�E�	y8�xt��g���,�1ϻ4ZL�7:����q�7���<U���·�ʪ���y�z1��Ae Ѻu9��%��8n=s?fy-|Da5G_J�8�t�ك��pK�7�Q}3K���p|g[	�Zq��Z��}rw�q�����9�T"д�OA|'���§wπˎ�$�߻�(�9A���h�IZr�'����Y'J�yMe���lu��ғ��g�*��o 'F�?6�������l�=�����<Js`�Òk��f��ն��~!�z�|�n���:�3-��=s!�E=7�՚g��h�{�hz�+��s���anP@k��D�#$>��ɟ&��1�5K	9p�3v:��ܩ.��,J�0T�����(M\��#b3���b��W�d���.�X���W��ל�f7�~�	��"�����{�����8#*
���Q!��5��jv�YafP;���mu�5	b�6J�ޠ�*�wLA Ƽ���~C>����BJd{�}Y�=OL>5xL�қ������PS��˜C��i��0sn0b�H��y����]ɟ��ҳ�S��F#:���#�ݘ�/���n�R��[��w0����y�/���O�����A+����zn#/�ب��-��#��q@ }.5���+/��_���?8�5~�n��󊱼�y�߫56=>cd5(ii�1�b�7��~��?���W�8�Qo ��}8�H|�'���I=
�豲���($M�=����F�r���n�n*�kK-���6�oǼJP���a��[����[���!��'�/Do���5�R�K���G���4�,mU.%��"�#fW&�ؕ�������m��a�T^��<^U��ֹCZ�_4��K��YT�;t��m2�?By*i A(�[Z��۶Lʬm:il>t	��HX�}�?Tu~rq���yf�]ݶ��~���mN6���p���B���q�\<����5�����kj��Sj�M뺦�&�1�S����Ck�� O�I�����T
�~��0��4Xu%�O^�2�]V\b��z�,͆�i���	��7��ȊX=m��eM��
aaE���9M@��.��M`Yv��������y��{>�X^���~Uͼ��$�6FZ�9y�<ۈ
'Z�b(��OO\�f�MXiR��l_����]Z���{��-�I�����W��0�c�S��І�ʛ����� u�Y������BUz�=_�Y5Fx�f?�����?�Y������t6��nys�����F���sPL�v-���Z�@����JcZ�>'.����з�J��B�t���76ú���v&� ���
x��<E��t�@���z�_<˷+帴���]`܄ X|�x^�B��aQ���Ǭ�u�~�0��A>����4�=��׏�b�VV���y]\�Ng	J�[�'K��� �-���m1'�����y�)^���V��ˣ��ycP����f4Cִw����a���ο25�����}�Bv"��ݶU5$�	�G�������!�#�aK[�]����(�-�f�J���T�+\����EN�tu-Q`N���5�'�N7���}�.�}5�ƛal�B��h�쑁E �i���޴��f�y�ڶd>��.�,��vj]� ����W�����*���M?޻LusgQsf���[�K"�c���=�;x�;1��=�}t6\�=�\^[��/�����+�|<)��P?Zu�z��cO�#�ۙ�A������?U��s7� L��i��1M���tk}�8��I¶���X�9
���s���5��qHė|7.G��*H/������  �k�깒賈a�F�	i%�����c=2�?Z��'��qW�У)�� �x�1�{7�ׅڀ�D_�����NEq��x�8/G��/�,�3���k �cW�Ty��������ccFMi6���eŅU�N��eSݾ�>�EY	�J��T�K�w[-lo?�ޜ|�+�xzsw��X���^R��Te&�6��. �a�\��n�I�K���I�,veS�?y"B�١<u�������o��+��^B�W7�'�>�~��c��܏����S;�������n�!���:^�kS�hϪ�в��$���� >s�9�\��Dމ"
Lv��
�:��{H�ډ"��&�,�En��/�Ӌ���;���R�����ӥ�|*����ғn��>�(�h���yе�p�3{"خ�>(�}R�D��{��M�ns��9�uZ)��ۻ6�65���(�˧9>�D���RI��3�57����햃�B�s[~D-Z��Q<�^d��j�=I�X~&��V�4���t�κ�0�z�]�Cǥ��D矝�Wz���v�G8Ŏk�]Иa����q�o?B�mf�!�2�;��i'�>֏+��l'�(�q1'�>ѿ���ZH��!k_$B���ڃ���|�d�wzl,YUC���c4��,I�A��?�}Z=3���IY��H�r�r"�*ȴ�~��d�v	��h��ܜ��`�.c�������o�����mw��S-��EhM��+���\�$ca�t���>-���\��ee	���]v<�[k�`�G�� ђvC��D���a������]+G�L>���6q�#�����~����Q���=c8�׀��i�a5j���~/��󚫣Њ�,�,��*�և2����>�Y*�.��8I�>�lC��@��/�e,-h~��ZZR�a3zB�׷+�(cm���p�U��;���9���*��y�%x�Ĺ�>�B����Wu��
���^�� �PtTD��nG�d���x�LHH��\`*x�[�ɦ���?��꜋�?���儰�g*Q��<�M��|������n��W���s4)��U�0f��c����o?X�[����d����q|���'��8��������03�+�7��T���
&E^R*W�����9b"^)l�ؖ�b��?P K���z�C�Pz)	ksS�[��M�\2�P���'9�!�Gix�Һ�PK���Ѳ�2��/�e�j��5�^���D��g����'��j�P�6;��l�ZZ�Ex�H�w�^x�L�*HؙO^tP���x�P��Aitj�-�iV���c� f9ָbEV>�Fɍ�+��.�c~C�NL�D|��i偳��/0,�zڝ}�.x<�1D�q��0�UUU�穁���q�,q\���@(w[��{2 )���&9/�P*e�9G��b�
?ɡ�V�0�f��--p��S'���W�mٷ�ڑ�P�DK���`��P�C��~M����n�gn�y�"qvX}{��k���nnw� ��.�m�FU�q��-:#��	�f�g�4p��*%�^O� j�9�h��?ߩ���y{����+Y�`v݉eLB�&k�@���״�������#Au�<5�f�]��^L-;�]f�2�wRynW� !ִ��^�}	2BB K�*^��3��;��e�G��mwq�Uk��� 7'�Y�#���<�ݪ�rYY�õ�-3cM�� �������z�i�h���-}z�ɽ�+rҕ��XTܮ��}��u��x�~�`��5w!X��U��~n�j�ZH�$o����Lr	kZ�*/�y/��A����A��C����'7�
�E��r���c,Rp&�Ut����@�v����>��ǲr��c;��'��(�7�U���Ը5: _Jt�K�����F����թ�5ZB�[��k��\ǭT��Y��쾙�}W�AX�!�"�'8�O����Xmv=�������b�����q5��D���@�0鏾t*�,�ua�����Zp�[�K�,G���� hq�&B�oUe�쇏b���89�W�\��A�o���m<u<<�=�.S�(�ۈ(	q�$���'��(t�z��pN�3���\��:[�I�j�R�4���0�7���k_4�U١CYiuD�Ղ��z
>�1l����?��-V��=F�Z�H�����z����L-	k���S~v�Gcn;T���7�s�q�I��Y����j��WT ����q�]B���1177��Y>���D~����g���6����d	['
`��3�����1�l7�'�*z���4�"�)��=�]Ȯ��3����bt� �O���s8�wQ�&���B0#�[E�l�`��Ǻ���m�S�	y�h�wHJ�I�I�l����Or�NQ�(��[R���"r� s�N�T}���ir!�a��Аl��s���!m�/�u��g�g]Wu=�!�; �r�Fz��͇�R���ւ{z4�z���4 ��VE�Uh��*-��� 0�C�O�I���2ǣ��������JN�w�QX%ʻo2E�>CHR�&�wn��l�IڀKCI���!,u�o�r��#�Ԩ6ɩ����ǯ{ο�7��#	���v^ty 钕��0}�%D�ݹx%uyo�zG��'�����?�����6<X`-�G]r=�H��f�/$#"B�m.�A�<iii)�
�x�>޲�����X
B�dB��S�>f�8�Q_P�T}�B��{�r����[��o�6B��2��b��rr������R�NGRS���S|��];Vn� &�'$]�8:�;�fw��9�M��3�/}��Z�z��i�����'D����(�C+6z�9���@�(s���Xb��?�'����zmc�*�P�I>g��/��99��/(
h����0I��7�Y�;F쭓~�ϗB-(*p�s�T2�L�Iۡ��&��n�D*b�>�>���a�*>���D
E�U����~8��"����[����(�":{���1���{L��*m��X%�px�q���i��o��"
�cza�~�(���	  B�*��-��^�=��^q�o��7
�G}������ܽ��4��L��4���%�,��Y0��i����R�d�g���-	a�]�S�j�K��7�(���J�"��ɟ�>���z��w�
~�y��..^��,��DA���e���AB��a�x.D��A��vP�C���c=�$y��[7�e���	�롴������v�dd"�9"6���2���5���r��I���6 ��>�U�j�$L��=_�w��1_�L��x��YȣW�΋���q�#������}՚+��W����
,����{�y^�.	^�����>�/4DZI�r���e��gj��������Θd�	�t� ]�Kb�хI�Z.I��1��0ځ$�} ���Ā^׵C��a��� �{}�ߵ����l�ٯ̓4�+!*9Z�Ɂ�Q�NK�����ү��F
�#h#("�S�O�ko��YK}��b��y�t�\ۉ:=��Ca��K��0�2�*��|���\~JH���ʚ�&H->~K�'-Y�=(���OQA��!
�`�/� d�Yי�̭�"o���J\�_� �!���{7��o5;��zd"z�P�^��v�-XL�(l�Fcj��1���!!KTҤ\�d>���3�SP7��P���	}>�P���& �ߛ��B�t���Xo����n��ɇ���i�9�7���R���y'K��k�����9�	��j�����2��4���2ώ�p�ܲ��5����ʹRpB\^����l��f�F��N��*���>�
$���qY�W,������2Y5d�e/��+�f��n�� �13v�O.�l(��Y���'�����`;!��v�~���S��g�f���|*�8A�c������_�2JDc�͆�������"X��!�o��vb���ѝP�WP�n!�L��?��qCʔ��$y��ǵ�ۑ���/@��ګA^	27$/���m��(߇�t<�h���We[���s-����q���***��,+"b�s����5��u�Sܔ�����j�;{\�ex�~P��9y$Aә�=8=��	����,D�),��qzگ�
���������ʿܦO�ka0�6�ǉ�ʼ�<N;=�O�}vQgE
g�͏��
�k����:ߩ$tTw���Ѓ]�B�^�ƃ����ח�?������jc��9�8��f�I����u� B��d���*���٣�s⻺��[:^��*=�˼y�!p����zF�vޛ� 	����C�}O}`��C���a|ś��婯���p7�C����J��I��ہ���Z����܉tK,~>+�c-�Z���#F3��Nq?��<,JU���Ԫ�lw�w*�=G\
%����7�5�iS6vv����Q�0h���'h�����
��z�j��Y m`9q9������b�(�$ `S;��Ӏ�$-��>4���ݝ���@$�[�-��C�\����VC���-��Χ<�����7�|�E"��Hز���99:��u��B�2gO�D���us���#���
T��.��U�X!����
O
�e���
��RC������������r�o"�g>��ԛQ�~���F��X�6s����/�{Z�33��0E���g�.*��#�&���$@a}��,�����+9��Z�T���jʞ�H_�<t�~���RY�I,~��e��M��D{}�҆EBK�����S�N��T�l�+�X�	��������		���q^͞�/گ��bB�D%)D�M �a����x������A���4�7MA@�ī�G������fu��iۖ	��]""44hw��A�E��j��,dhHT6>��O��T�z3jdo:w�{�Q�/��L!����b�}�r���������h�@D��C2��N�����@�X�I.S��Đ�%*��sD����X&]h��ȳ$&��l�~�p��ԧ�c��2���)1��6lD�}馋��J�6o���I�V��`���٧�]U`�W1�J-֠h\���̓8�\�,i���R�E�����ô^EOu��3�	7-6z��In�4M�"�
�.�4]R :�����Dv�������eM�q�0�A д�sɊ�Ռ��" ���?d"�PWȚ.%�����=��OG��T��^�B�y���Wf����ن�D�<uBB)��!��&_S�W��h���Y2�w����C-�訠UN�Eӹ1���%�,ߔ��ڭ���V(,�/{,p�ZA6�;D6�V�X�v,��  7��|L��<0�tBV�w�ɲ̐w�-�aT��vw�F��q����G���63�Te��"~`B���Ԙ;?3�_��[�`��>f��!��.j����&&D[D����l�NY�Z��\\�xa���n#RA�U��É+x~��\M
��&�<�T������g8睿�s	/ M�+4@��|o`P~��}⯙�����F�:F㹊����O�cWA#�?�<.�'���\�թ����UH�0ek�[E����\%y��-����I��m'�gm�b�F���D��e;���*+=<�?EHr������������\���Vf�x����m�i���=��˘���3�[��pp�[+%���D'���v�+�ǝ#�+UB2���M�0 �̝��b��P!A�0KH��Jc��o��Cr*�2�%d���g�[�F&f{��+����~#��L0�|Keg�^�Y���d���T��Bk+����ԧ��Xk�"�^BA���C�k՛u)c$�Q%��!���7�cE��*ʾ���o ���
ԁ�ځ��Y���L�Q��5_y���H�#�̻�u%�J����@�*/�R�R�����nntw�����b��I./&,��ǆ]>zdd�_%:$םa쐮-R��Mj�� ��2�/������Z�I?K���r�zh��?�|�RҊU,wI�Ӌ�?%.��è�(�!�,,v��f��	
n`ȉ����X��l��t��	��ּ�\K�A��_hםe4�e"����ޥoj
%��U�avV���1�P_b ���Id�:sBa�s*���+ܦ��.���L�;��<�Xr;"�/Ύ��~��c���7\q���B��z�Lu{��u�#�Ȼ#��d\�*.�u���䯒��4Kj��2	@TDY�ʬ����)�l�ԽC�:yڡG�����X��1l���~
�%u�Yg�+	�s@[W��ә���fMٮK���
�o����?&"�k;�n��9�B[Y k�N�k���������e�6���Jq�/�\.JnD�"��yt���1�e� Hw%}�;,d��@,���4�3����r����?*z�z �{-�B��FBC�9nh�� t�?!�����*�{�
_�N��/e���>�n�`�ͺ8�4,�8�4A�b��÷�I�A�'O��qg��櫪nx���ų�P���	���Qm��隴�b���,C����{�>�� [�L5t���-Z���&�Sd)g<Ā ʐ��PDQ@κjUe�<:��dFl.���by�%(���nGKKU�zqbGdg��bWۍ��i�#ԂQl�����i��$dee������JGF�a����c�-Iu��V<_1y�&��HC�O/�^H��s�3�V��8'9��&��CM�O!��_6;5 �'��X3J��+���{6!,>?��l��9Oprr�J*���(0�>��jB�<��ʉ�d���bL�v�`T�_Fbak��)���{�/$@�s�WJ1U���٧����W���
(���ؗ�ׇ��ř0�9�x
Ԙ�jc��-���I似xr���k�������k_0sh�h(�4i�ǮR~�
��~�(Y��� �f
�d���Y���*��d������deF߁*�� �z��� �a��c����u�	^��O��|��.�x�L x�9�ז�*�9A�9!s��%����܈gZ���@7�%��r'���T��[������zWJ�K/<��ˉ�~k��Q6�������j%�vd4��e^�-�i�g��@��A����7�л%4���P��ͯ�������&Y���G��)����(]�����n�K2?h$�����O������G��\�&&��U�y F[O�U������f����b�����l���͖��̞�zQ�	H ���LI�Ҁe�N�JHԵ�F������h}���|l4_E4I\PP@=��zvs�<��N�_���+.�zC?
���W�|yt͌GGW�J��C���>�\������-��~�ej!�w#�#+Y&/��B'�M����E�^�/!�M%3�\��#aH	�	�����-��-�k�wW_ +����1z�;�r���!�w�����j4Mbb���?J��]��P
W�&�$�� ��Y0�z�Y��܃=IkQ�X�NO����6���ʂ�!��?Xg�X�����Hgrb���h�=�d<�e����{ɧ�Ut?�dͪ�@A��Z��K�����/�99�2H��/+c�T� 2���x����26t�="ڧz�����~K�R�[ZaȘA*P��b���2��{L��N�Q�L�lPA����3�u�Uw`l0�wi��"P+f����P�_^\�ʗB������Ip_4�8�����G�y �xC����!�$UE[�}sK2�/��3�*<DdRoUk��D������ �����#W~�h@�9[�����0R8|B�5�p����&D��lS4��c_��|}]��B��3�J����N8f�ma2��r����8�Ϫ�����F�]�#��2�XQ�~���`Ԅm��E���!����7w�W��{�k�͸��!�������*]f�{}� z6p��:�|PQǂ�����Ժe���MK��h�3�qC�%q�����J��lYJ5��d$~�H ��}"`� ������L��\=�؉�-�8(�g%o�c�P�㭖�"��+]��C�N4(�oT��iVP_d<�>J>���[�As�r��!h���'X/�J1��_9L�W>8��8?���˯��^ޜ��N�B��v�7���V�^� G�L�)�ǆ��q�!��K�	��IA#os�{���<.�t����:))z�f\_nkP���"�(|����Η ����iX�Kǜ�Q�� d����Ū�Pƽ���9�)&��m�s}�V.��^���
x����@���[�&s����/Ɣ�W����]��U���5��ʝ!z���V@k�څ��c0cښ�G��뼿���G"���Z'?��Q���oή�Vz2�� ��\��U�t^�r|87o9}���VQ@5+4p�Hp���a/v�Y�Ɉ.� ����nY�؜��ƓV��������6�,M�H+)�9v������Sʴm�O�@Q"��+5�2�C*���������@8���C,Z�/.�)�²nO�Iﶵ�S����r7ͧx�(U��he��?\s�v�*'�T'feEѩ�赻*T�`a崴�W����?K��58��@΄��K��Ӕ*�<���FW�2$�&����V�)	�.����3iC�K�-���q?hN������|�HV�:��+<X88܋�Y��~uuu����-�+M�����=Z`Ei�@�_��2����c�,�K�X�J4��*��� �5�y6�P���nH�t>!��\�(K��ϗ����+F6���MJG��pu?����9�T����Qi8-�)���
h���̴n�w	ߤ	N�D 5 Da���5dhIc̲]�L���ߺ���J�
�� ��݌7��S_ƭ��
޺�B }�Ωծw�v*�E�uCAN>��q�X���`�6���R��_����ߠ��O�BN� ����ƆN�[��g�ˍb��@���Ы�2�t+�p/���=��%����B����=nB�=<���̨���5�����"-(��^nb���]rM�`��Iȗa.� �����E�����1�g	5��s�Ug:GH.�zB&�a�7�Br����)��2���{C=�11�{JE��m�E�=�F��F`�~2�f�g�T�tT�b�~������������U�A��s������ֈfuQ������C���7���֠�o�o)�0�G��$�D���U�3� ���U�y�׺��q?�ZVK�@wZ�L���B1i� i�P����SQ�ĕ��L>Z�����V^��cC�~|m��$>�>����2>9$`�%�s=N��~{-!�����W"���[c��+�^�Q�/Y��׀�ݛ�w8(-�5a��WRT�tw�EU��n���p�����#��@�!4�\�����!n$~s��ۀGY���- ��L�؆�����te���/B��la{��>�oų�i��E�EQ����SA��'H�5�(��I �F �y�v=2�\}K�#�E��]���:�J����3oxnJ�n�=�e����I�E����]�r����������g5_����@)3E�x���وd�=?}�<�E��[�IM�{����{L��-����eh �lv��q�ϡ��%�[���֫F= ���e�d�Ӷ�����ʿ����TEC����.M'��:3$D�f5F���'�j!%з��mM�9ˊo�e3��'���A_Ƅ�����Vɳ�귔�����q�Ci��*��x~�AHsI[[f��#v�0(i�lA��>��%���b'�H��Â�%
B�R1���]�?K���)�dǗt�ޠGV �&��)|�!mA6C���!���TF���&�Ř���*���!wY����]BF��o�[)�#q����?ι��Һu�QN?�L�!������v�CuwY6�TN�g<��n]P�H�������E�R
�<IY� :��=\є�V>���T38�&��gG>k1%� iR�@�a�d(��^�&5@@��*��B	�e�.�t���V�8yv��U1���pY�H^���v��c�$���O׈��h��������d�2l��	�+x�U�ק>��V�8��f߆1��Y�8GPY�NB���E�I��:6�#��R���W�NMM�w�0IHLD^rr0�D�]���Ɂ��L]s�i������͉^3��g|Y��"�&21R��ڬ/�D~�VU�#�b�����ck�ħE�Z����N��c6�.�z:g* H�<���?��s����U���22��	��w�8��CR���<Ѻ�;8���F�(E^:뽾<1�$�8�߉��C�m�L�D�2�bQ�˝��w��R�h�������h�ڈ$Pa��"QMHJ2����0cK�Uo����-2eO�
v�Q��
h(�rϭ���`NƷ�}AU�Γ�n �IH���w��X"�)�a��c�G�C<�v�����d�t:�|P�\N���c
�����▇�����a��˨(P�u��3e mg>���Z���5�\�.��d��U��E�А���0P�DH��̪v]*�䲔���晥�!y߻U71%*�?�_�#��������#Rd��� �dccs���dԓչw:�Kx�x_У�Y�M���t�����0���	���y+�m\����,�P
˕´�?�U����x���٧y�SX�7�{M;24���1�9�X�k��UU{��׭�आ�0-�w ����d����_��G�`тON�9��$�6^�s&�.w��pT���'dDl�s̟Wj��"rY�W�[����ښ�f���r8�7� �}n^�b#^,h-uMC�g!����������Hn�y>_�
�Giq,���ua�)�|��S�ǥ�J�>7J��9Y�2�uKx��F�����n�����5��X
+.'H=����E�ֶ��,�3� ��~%��[KP�b�/�؅�77��"�q������>,'��X��4��s���H ��	�����U���6%�� ��b�=��nd�a��V���1I���[ɀ�u�L3#Xz��a����Q�,�**$@����A{�zi99FIg��
��-�-?x�b�2<7ư���frk]���Ѓoʓ> ���L���5�4sNOO�ZNQ^Σ�=up��W�	`���]Ɍ'���)<�@a��lCOdC������!.惏����B� o٠k��'��)�@Fq���Yzq�#���(�o~s:�	���L�7t
��@��y#�P`�|�j��]�C�����/����_|����A�X��M=�V��B&��rY� �~��B�ۿG̰�!�tǨ��6���ʤY�g�+
���D�ju�1â�1(����?]�_SSs����BDYYٴ1O�.������z��= ��ȷ��Rb���V�ƤH�Jk�����w:��y��fryHe���������H[<��iM�@�8�2�h19%�M�'G��|��(|}�o����N�GW���p�9�I�J������0�5)#>���x}�i�YI��ڎbfd��y�5��T������9�����С<Y�
� c
Q�/��ܝ<��G�%!�f999m��ulll�O�,uz����n$��hnl��/1���+�p0)�9�ׇ���GT_>����&w5U~������yD����]�<n�f�_{_����?T�B"B(�R��c+["K�([BvY����^�,S	1��c�(C���G����������^�>��5�3Ϲ�}���z��<���[ڛbNy)H�q7���vhg��L��NN�߬t����p�.��_�wD�:��j-n^Q������7�l�]�d��TVI��UX�="(r��D`cY\� ��
��G�W�DA����c��ݿ�� D����(�� _C������`��+���o�zѯ#]ëL>y�-��. ��"&��w[0���
�o�g𴇂��38��7�'�o�{���M5��=��j�YP�'���I�� 5|k����	q8~���U�##����楎��v����1|�_�&	
�˱˻5P�]T{���c*`�gW�ܾx�q���ل�D�P��CƐ �iLzD?�jsz凅���]Y�!�Z��g`a1��)��S�;w�Ɛ"p�Ѻ�X����3PG3�R)�9?BN뗘%�l��Do2���7/�q�������5�m���Y�ܽy���(Y�?7��U���V�#��NM֜�B+^���MC�����u���,W	j�l�]�n~!T;������Rt�D�˗^lɂdѾ��!X3�.�늘�b(\>��1xd��%bP�}���cEw��@�����X������Y ��ŝ�ΐ�`�Q�S54@?��oe�����h��m�B[-sO�rso�G!��n������[[^�'��G,����>�Dj�������0���
Eq�f��H�������L��A�|����>���=	"�|���������[��
��;�܊��r��=��˃��3@�b>w<y6���uɁ	����Ȼ��dl�B�Ĥ�����"�ٕnʩ���-9��l�G��h�����f����A�-�E�:����.f��L�S|�!k5�b��V�~Ŝ�u^R��^pd�@+8���l\(�v�º��Z�P:WO1A;ņRO%��_��J�q���:qF�����ݭ�WcÀ-��]d�e�~eB��KyR,���3��<}Vˇ��@R �}}*I�oZ�(��``��� xA�%���f�J׽+g�����h4����M�:x����ҋ��\��G��i߶��^d�>!i�������~��rY0�[�ͼ�#~�b�P��C5�����(���oQ~|#�qGe]5_�_��3ϸS��oO�t�~ݙ=^p8�1�eXpS(q[v*���~�ңRO��bF��@(��q�)�)��Jw�\ۮ){O:$ ���ҏ�Ykj}���j�������pj�oTaH��[:0�6OW�%;��]���0d����^��y��b�����"ۭB9�4���uqHe h&�s��I�2]�4h�U>�&�}��}#�QU�$Uj�{���n��iv��HSh��#�!<d>
�,Ӗ�=��������tˡT@V3]�pa��7�����Hd{;�+�}u�DXF�|�_����ǒ-���GN\��r;�Hb+5,^J����D���D9&*�������1�Q�'41$��Ͱ�ZLs/Q���;w�&Q��������_�U\72J���#���=]�M����WX!j�p�T��v!c\�������%��Z�wn���5G?�mi��}��$t�m�.�GDH������4w��w��6�����5�7���c~Z���:�$s�@���d8� M{fyX;��晡����JI�t���@FX��m͝��?%Ư9���#tdZS�|� �����Ҹ||���ś��$���騵g�1C�	tn��� ⍘��NP�T�xQK<�
��F7��0}|����c�'9�D20*Y��v͕+��-��i�o�Y�
��U�ɑRZ@��5
"h�稪�Ў����8.N����V.��7�;��c�1Yr��N��:���L	���p��9�uBV���E�̋��#�n��NCB�����ˡI��Zq�"�.5���2r˨���
�B���t��2V�k���=���23���߿I��?>Y��E����ԲxVˆ[��/?a/
5�Nt{vgO���@^#�̓���������mufĻ�E���<I&�Ύ�����7�t��H`FOO�b5�����vV�vV��� 2O��8I|�0�.�ՠX7ޛ��3�r�0�����cCA� 	#��ft��K����I9�����{Ɵ�6�d��E2}��U&�����/�͵j�?_L�O�����} l��j�6����ۧ���?��@�88��RK��0�����F�1OO��&{��o�]l �!�
�`N�b�ӎb5G��\<'>���g��UkHT�zA��1�����&�|��Eٌ;�pC�����/\�����R�/�v�-���,�R�,oo1K�R`�#P���]Q�w&0��
,<j<�7�* ���>u���-�&�����9��4"��-���6?b[mS�#���ۖ999���АEW(	_��<s�(��������Z^�u��ɧ=�}��d�ә;SI�{3:��Ѱ[F�z�~I{���_=�x�s��h����g��;�[��Re����H�5#�dч����M�	�o�,AmUt�A|JJ^�T��R�HC �8�.��q0l(z/(M�rO�\y��5&��X&ۿ�E��r�?�|ǐ
�4��ȕ���k�$v���P��ܠ�D(�C.��Ί�xg_n�d�~���C�3��z'm�������b����5���NQ�H =�C��s��f��:���0v�앾��N=��!����1(�XJS[���2Yq����׌�Y��!;2����v��4� R���ul��~�F�,Z����!�'z�%���"��@�E6
S@��?�~:���qΐ�����ŌR�h�����Z=�,����4o����}��#�H��~��Y��c��h��J7��K��b2BE�V����a�z��7���	^�ř�G�XG���	�Ꙡ��ϟ����˕)��|�"l�FOZhv)$�@Ba�s/~G�{h><-�����R��/���y��4p�2p���W�p+	�ґ7z�
��!�$3�m�A���x��_���� �Y�/���x7����S.M8]���>�=cip�*[ �i�p�i9Z�FW�5��/��V��=N�e���GBu���g�9)�k���,�u�O��;9??����"���Z²���=���<y�[�p�C����aw}XB��'�vY�)n�\���V�=1���t7]FS.$}r[���ԡ��w1�����2%��￉�e�����#_��b��z�qP�QNUé�1�54�
�~���ˇ������]M����h�Y�U������b_3����˘��A��'$#j?��	���6�u��ih)
�2tKXq�;��#z�.���?�UK���D�Ӄ��O(@�蔈�M��W'B(G �ؑ�3�g��>����`����o��a�POD��-`)iiPݾn��#��nTR���,�6+>9�bqc�L*~˶�u^T�8�ų���������a�gA�iM�O�;q�'�ď@+v�0H�|�Pd��+�>C�ĭ��H|\��[�q���
?p�+|�ՅR��<�iD�&����&���h-u���x��֛ЍI�<�����!���{�D�P���h�R���4�
��&CS��3�B
\2�$:#�����T�ϩ�M��KK��۩v�u6�)� ib��Te.�P��G2�_�[Q{��S���x<$��?�����x.�`T{�t�r����ײ��"��]�x�{��V�*��H�Ę�/��6/]�ї ��47~K���^Y���1��ɽwZ$��Y����Xm%���c�nZ��B���g2kؙ��ʐ��7L��eHJ��d{
*�{�?�e�3j".< 6��>s�N"��f�o��
L����7��uf����%��?��)��������A�����j-�q�a�K�<���AwP�-'�G�0Y?��ohbB�ahUn��������n������P��EЩɡ��P��>�I��U��d7�y)�d�L�����c5�j���ʖ6���**�`�c���ڇ��qA�n��Y^|�W��b�F3xr��.p'�ؕ~|P�*"*�&qF����Im��&�P���'��S���x����ٗ���[����#�0�oߪ�ݖ�j}t=E�*p�R����b��@5�LtlO-Q�K�λ�����\����&�����$�?�1v7c������Ɵ1�^�'�)��%�>�$[�t����>`(V޼<e)�����T��7l�Lv��VlV�m��'�D���F|rr��D��aF� =��y�:��ʈ�WF�$r2�r>����?�^�����?���|���No�e���G�>@Yc���ĎNN,LQ֕c	))Q++� QCN7������U�+�ru�X�,��*��V�W.�z��E�1���\�#�XŒ���Y��.^P��N/�8�p�3�N;)GGǓP�df���)�B̆!=��X�:���yu��_<�w�ށ�������-�5����9��O�?w�]n��r�|���|'�BcQc����@bB����1�0���J&=!--�LL��=S�׸��v�I�5����Q8���%ݏ>�KtV�gq?� �����h'���{L�w��֙����2F�s�Z���`o�ύ���306�C��Իv�Z�c��JJ<�4�q8�!x��5aC�$V&�L�>����vS�oڌ�����j�f4oC�۷/���o�)�E6��{t �X�_�,#�ǡp���poɺ�,�ŒI����a�0�<V�ϟS
��;מ�����&���`4����)���T�S0���Y���s����]�m9Y�3��c!��ov8z���PP��R��.C�[�n1�o-��^>�Z���h�
 B�޽a����`ur�����t.���OE_�gT`�6L�Zl�7���
6�ď�x��2��_�%��N��n�Y�������"�z
���x-P��F]~�@<D}����C!���4�#Z0&��K^�R�\~�� ���4|,V�<�P��q��_��ץ��QvR���㫝�@�mlx�91�Vr322� �`'�ڃ&�<�����]�`�[�;�������2 �_2;x�ԏ�*.�2���=!�^W<��(�e������q�h֜'�m��Z�#�Zg=�K��(������Q����M���.�Կ��H���[O�b4+**z���[���'0�h��;�x��`��n����L�� ���mr@^_����=#���K�?�q�P�|."�-���Z!�~��������<(��ߔB��hol���H8�~^�9��.�Ծ{�7G���^�jc�1��p��reM2�����'s��y/,�������`
ބO>P.B1�b�ӄ5�ia��\|�Or�ۅ�T�?�H��0F�(��yue)������x�IJ2����T��U��8��p�?�K<�sqk�|�K��޾�:�{��p�8nq�׬l�T�'F>zPj_�G'b)zHxq"�?x4!@���H�c�&o���Z㑑�џ?�Qy�2R��)�Zqv��b�MS����ʎڼ�+s:)���9��#?��Y�p��%�<�w�����W�Gh��R��6�����`�}G}a��G�eoW	���=�wѴx}�W�9���4�j���Z�I����>���Ƣ�_���s,7SȌU3Sr�6�+I���-�|��3/%}��^��Xhs���6+4~��KNNv�ep��1���3M�J��dA�#T�qh��`�����s��|�����V�p`yXp�"�jTJ�f�k�y|�H@=;�;N����񠞴��i��]�k��z�is�N8��ᢥ�Y���i\-���M�x�1�����1B�7���M�G�ʖ{�yn����b�W�M�sR�T�O�����������d���.��q�x����nF�r��ڴb�^�wC�f[t�r̈́��E]�'����f�N�s�g�[iҏ����{�vnM�<��<�ő�����!��ݳ[�2���2r���&����7��/(>�Hc�ͻ��[�Y�fYU|�V�ȵ_gC6�U��+����X�n�^������Wg��(�s{-�k���7�1���?~"x��e嫮�{s�>�T>s_��<y�Veؓ6�����<���$����*/��_�jl8_u�v�4͜w���]�QA�O�R�����9�.��'R����0�t�M�8�-:#�s������:Q�|wO��������.9�4h���H(ľ�q�YN�?^����t��#�C���"nnãa7
���P��z?��Л]e�����=�|�4�2y\|n��Ӏ�_0�N j����}b2C���>�
���� '�x������͎�Ŋ��^��jK��x����:c.{���OQ�\g�0^���;�m����� �8���+m���V.�5�4�C��T�Ⴌ�G��aT��~dw���Ĉ�$�W/*>�&�ߔ߬�����{as2�y� ��ss��./?;2�2[��7HWy}��VLQQ�B+�e�|�=��3�<�̟�����9ԡ��uh���*m!�@�Bԁ����r~n�$�g{_�2�!U�����d�����d�	�ZX�w<a:�|~ߟ7L&FG/�؂9lÝ��l# �6]�����:j�G�J��d��yQK����N��Ok�Z��zgw���LN�3E�vp�G�l� em�Wxz>*�Bvw�?�/��}�rx.����R��.ܓ
y:�nJ�^����ё9T��b��-�=���Xt99�E�Ȅ(o%�m����U��u�6q�{�(lD���L]�O�o�+iŞ�����s,������:�ܪ��`����Dc૝�fW0��QK��{}Ŭ��';6�ڑ�	l}��Zc�G��|*�&�Y�?��p.��x��A6�t����Gi�Gd=u�V�p�S�[̖����A�:99�����]M�|��?-3o���#vv�;wi��[S6v�z�2�Z��tm(�������92v��I<������(�iF: O}G,߯a���u��3�9:)%���V����٤�$?����L���l����:Q3�֦)fِ�ݯ(�M��(g�����i�鿶��7˃U�,/��:N���{AI]��Xg6AKr��e�+B�+�c����}B�R��f�l%�|6.���$���\�r���[�eڽS��$�,1��bc�N�obe����*�L�r�..�Y%^*O/g�����������m@ �p���C��.z�?��?��p��A&C����:����l�I��&��Qz&��?�"�R!�&���ŶwQBl,F��פT�T�Ȭ�E�� =@��K���ډ����y�P¶��C�5���mŒ��Z2p�/}^!���-fWP�~Z�O�9uJK5�\LR�eo[�� e������Z	���`�"��d�\�|��f��1��ܙ�?|8���hl7�/!!�������VAe��EΪ�k阳
^"���<������(��1�O ��.��J���tX7H�`/QR�\��C�����G��o���H�k޷��d<�u~o��U���b�[H[Q�����
0uq�	���KK�K��vvv�	_{''�q�. 4�SR�l�B�Q�����i�ζ777K{6��|pM%mow�P¨:����g}�\٫	��J1Ⅾ�WY�>X�=w/7�}�F���ؘ��9���[@;�k���t����EEE��jօƢǏ7��&~�M��9���4��	�	�B��!g�ݵ鲱պ�Q'�3� i"L~˧��d?00Ѓ�����w�ƕ�@�i�hf_\[q�����֧�UV}������K� {��hqP�N��,FW}�H."�;�з*�N���2[�0E����@�n���t���>� ��E�\��9�?>�p��RR�R|�&2�J!���p��|h9����pm��r�B3���6(H)��J� �;{�1ff��f��U)Ga�F Qa;�4���f�2	��`. �iB��uE#�E({))�l�K���Xu,��N\��)�9�C�����TT$[�d�޵�Y
N N������Ya��@�g��k-��C@p�^ ���ǧ��!��8���NFq�|���/"�k���)�i:֌��j�����z�G�����i%�쐑��t�=i��-$,<�	�j�حŗ�l��� .���/z�;!W��E"���{�vę�s,Py���A�����1k���B��,�!22:��[XXФ-Ү�i%��%����peee|%�3\:���[�YZV� �&?A��>�߮u�;�}rM߯0<?���6�jpvs�6�<>Tb��x��ݻ�fCu!�&�0X�X;�C�����V��&���l%q�r�6���58h�P-�ǫ�@t���8�����:�#�,���APC���![��W�+�
M�ژ�Z���|���/ �V/���h���yߐ�M/p��ʤ�$�����]ͯ�Lc(\��Q׷�rnmx��`�9��z��5�8T0�̉I��&+w��{fFF � �4	ͭ���Q:������
U����j�w2B*�|�4{6��| ���%G]�p\!��:��@	w��h6 29�/Gz�vQ���K���i�zx��SD��}�I(����Qu��_�����������q̊��[G|�{�a�ecW��9t0^��n�����Zc���$ѴLcL�`�� ;�����6V���bLOh<�y������{`�A��������ެ�*}��t�u%\
�5�j����!�cxkKş�}���V;� ��j��-�A���W۹�#��7P���RcE}w�A�5�ԋnX=�?PK   <?Xv����' dX /   images/afde01cf-9dc8-4de2-b588-5b54baed9cea.png�y8�m�<R)�R��,I%�RH���nK��E��"e/���NY�2ɾoe�ؗ��f��������s�5����s~��;�<��P�C�F��`��^R���l��`�����Ի>E���|AUw���a ���x���9\��G��JW><�|�E�ᶋ�w-0nnn'��m���s�8�p�2�$Æ���*��u�����J��\^,L�}��tc[Б#��	��ި���E�4��ź�Z7��~5�kͻ�g^-YS�2�o�]���;g�+��i_�ʒ���j �&����t��(�+<wC��a�)d����KLMI\�j�Fተa���[����,��Ν�U��_���pp��k	wh�:S��\�A�dP�$S�dC��G�Czv��B�sc�QԦ2SZ�I��y�t��jem-U��E�!��/Ot(9�S���!跴��v67�}�%�ygF��y���j'	��&�5������ҷ�WxL��T��T��"���^�6�5�$jc0��@G��b����Ly<C�LN�!I�a%���K*K����V̳(CFLH� C�Q�߭���JՏZp�߈s�X,?~�8>�k��3��3���0��VK[�ۓXE*rǳy����_�ӎ�
����=�<_!D>���8QD���Uq�^�p��Ymm-A���{(���� ��7�Eq�Z�0��é==X�K`s@�����������(���>��q_��L��J�-�]�ݎp,"3��
�;H%g繜�Y�����sd�k�=6BGc��Dr�tBi0���e���hRa��a�xddDl�T�~����B�!
��m��:y=�S��4�)	�\v�K�֔%��C����tt�n��3M*�}|:-+�awc*3z�ʃ �DMl�e!˦���$7q!�@I���3Av�K��j�	'����G������DO�#��-:�aq,vs&
c&�&^F2�*�Ӷ�*�l������PY�2��4��Z�/L9�Ӳ��8�����7��Իp�(����5��0�o�>-���3��h�P��k�'c��H+�7�5��2'�i��[�,颬����d�hܪ�(F��4�;
�	ou���%7V&WC�.��pq��ks��佘7Rxr�SPX|oM���v=�}��-����O6�2���9�f]�"Ʒ~�M���,ƘO��<%�뢩I�er�G.͜���ݥ�IY��<!nm������v��R��2��ţf�뿬Rb�w�d�ǆ�oj!zo���c����Z��S��B�F�^؁�����ˤ���ѷ���T	��r����?I��_���$��Jx�0o<��ap�V�����g-p2}��H������y̍�%�m�����`����|sAظ��4n�Q�z&�б�O��˳�����Cm����l��o(~��Z�ʽJ��7����o��1���8N�*<���C#@����|_J��_�߿�t#rb��e��6�Ta�׶Hi7�u�:������]5/-:ۣ��壱t�g!��X(Uk(m����|�9�w}�U͙fz���w]e����bH��nQ_������B��&%�s���͐�=�:�pλy������f�h����������;�T&��((�Ի啴�E�k���v����?]^�6-�!�Ed�Ppz1���˳��Lq��f�B�������Ѷup���5��}Q��E�o�>
72�H�@1�Y�A�K=X1D�o-�A+�-�D�w9{����3�8W|��`X�C'hty+rh��6��������饣�,�����n��Cʜ�o�ь�]�|���x{�!�}Nf�&u���1J,�JW_q��I�Vb�����a/�WK��v
(D@:���T�âƐ���'�F.�8�����3��z�{h꿔ẕ��l^$r�'1���mX�(����# *W=��9έ�Y�0�\!bR������3�6l����>�ja����նZ��0yf`��,��s�yy}��6��|�j��*C� Pe��#?�G\;@m�թ7ܻ�$��]��[P����\yur���ڥ��Og�~7�b�,�#q�^����#g��/G�����H��"�y
rR�� ó��L�<d���K�����l�3�|6?�[�S/�E�4�:!�U`�0��O{�㝦3p�.�S7�G��#V���z(�c- �����"ge�'i�)�� ��t�$�!��/�B���pd�%G�K����sD�.��fn�����0��	��`��+++�JJf �@��m\�%�Hc|��Nh�F" ������͝��}���1dz|ʍԳ�ng�5�N��`������ �u�A%Hȑ�k�2b0��*ϑ��
FF��p|zL���;�T0�	mst<7����~%n�U2\Z����v��i�5�]���z2o�X��O �����^��E��|��AL8M�a^T�{t�&&'c㰴z�A��nk��e`�T�KH�4{h�a:�L6��)4h/��ܴ4q�ص�-��k�jiKE۴A!���<��D��c0���?C��r��ά����G�a/FA,���i<�v}u1T��~�H�)̥/`����?�H�M�SЛ��jK�FqUp�S4�ր-�\�lS�������ؐ�*����w܉{0Z�A�p�rҋ��Lw�W��e���W	�D�{2��B�j_�D������ƑH�[(Ԁֻ�ɩ��z��H�Y�gX��L-�%��p=?B�e����u�jqkk�����5<��?ҾjLފ���O��q-�in8]QH� �������x�/7tl��7;����b��TqR�������\r璬o��� 	����=��O(�3��>( B%��I�4�TWZ��mf@����72�itZ�6
�	*J�'���>�'�0�
�D;����:X��5��Uq�Pć��i(� �k�"%|���2�ؼ�`@�jx��%���=��Ŗ����cJ}����
���WZn��@=u%b��l�bבZ����ԓO�i��$v�1���)?�Gi�c���4�W�+��Ց��/�c��Q������ܓ�W�o�]Me;I��T����*�R��2PZ����Q�3V޺X�GUƂ�7�рq'��T8xo��+����.َp���/�H=!�Ws̖��+�T��_�] �HU�ݿB����S�Z���[g�
�c��}T�G.�d�x�[�J�mg�m�0��>� Y�9��S�:�J�E��i�*�A�T�{'�"E����mCu4F傋���S?#U�ӰoO�_Y�{{|�B�����Ž�{L�W����g}�T=ބ+-*m],��u�ES�qJ��ՏWJ�r��{�B.�w�R|��f���Sϕ+T����m]��D��.w���lԃ�B����	���6r̘����A�{{�(8��JI=��{��T�d��v䯒�$�cx����^�{��Tt���'$�#x����Ǽ÷.�8Q�@f�}0པ���U�}=�ףT�[5]�<X}[���{$UG������p����)R�^��]��\�U�rLL�����Ww��zaVzUI������Y������������e���-H�c �	iJAכ��?{���o�����'��
5�U�	�;�Q}Zٴ��D{���g�\˽;(�a���$�2koS�y�d-U�n�������P����y����W��>\����x�	�*D�?#m�x�
3��p @�Vʖ�j.�'��{���T����'-�t�b}GV�y��z*�ֻI�[N�3��2�*��w�7��G���o&�٧k���lݸ���ֽ=5T���5������t�b���D��Ԩ,^��O9ml���?Q����{��|��fs'�x���zO��Kv�?�-qB�r���yLU�����=�'�$7`閮���⿥ZLMe1���̨�+~�?���rCH���ӧ�yq��a���q��;��T�I�)-�$i��v��l�=(�������=l,�+d�dv@ �v%//��C�������ƈħ$�}�86P�[�����B�W-����y��<{Ir�[N����@����0ӥ�AQ�ꀃr��dB�7��/P��j]��yE��1V�l�1���퀴)h���U!>ѭ�jL�5Tc?�t�?�R��o�JhHS�J���gJ�TՒ{�O��#�����p���3�_qX�V^�C���	��r�A���k�w2�^�6��6�9�q/n����?E���9�>����4K��u!����9��׌��I���Wnv�F�mI��9ێ�6m���V]`�}U3�.o �D���Й�jj�r���l<*!j��߇�c5�]������b�wJ����Ǌ]!��B����7��-��s�Ź�%��clڳ���;g��_"S�h����c
<Y���k&p�U��\����x���n|�_���e�����3�̌us�J�	:t�te~�)ۤ�řR4f���9�5O��f�̾G����\�!)�B�f]��~�ԯo�(=nK��P��C_)�4\y�6mT+n�X�+)������Z���+f#�"Em;>P�nA����Zk*{��mJC�Vgv̸	:�,Z��\�)_,acg�+���ͭnmyn�U�Z�h��m�`R=d�é[����ن�􌬧�i��(]sOG����M���ر�w4A�v��S$%���ǔ=�\K
��H5k-}}}��/<3&��g�<�Tp9���6�գX�,	!ډ��( �f�G�p�3C5�G=�����ǌ����LL(~��d���"_`�)UX��mJ�)�q�mѹ���Tv�o�<��o�wӵU���@
��߂���n��qm7jjm}�e��/\��n�~��yHdcHd�]��e�mh9C���*~�Qڬ3�"-��5�ܺv��n��fff�k�\��޳a��_�Q�0���s������A��U�֮���t<�8%!ɟ�/w�Lq����a���Z��d�����]h��eK���Lk��d7$g��Zm�E�Iܞ���@����r�E=
 �U��8m,��9�q�BJ�������/.r25y�7y��=좦J��&!WN���*%��	��B������������A�Mq:���l�,�L�YՇ��y��ɫ!3SݢC��w�w����]�?}e�q>�-�c8�^F>�@C�k1�k�y���)qT����u�����ܷ3��, ́�|�=�vT~s%��)�I���kQ���:bk�̝i�?
��.C�ڴ �ۘ�ހ��(�m�D\�#���y-tRS���K�z/`�qbm'��jW; *SZ
��ܱ��%Rzꆡ���%��R��-ȣlm���+�����ٳ�(Ȩ�G���)�c��64(|��|8ڍ܌Ξ]zK��0��6&����j�13�`�kO�����Wu|��_S32�P���o<%�����OZ3�S�.�c��6F(�1Ȼ]�3��!��&�A���Bd:�ݵ ���,&e3�+^��̵�H<Di}�Q�y. �*ō��������
^S�gC��wm���򯃐1B&�2d��6��$�������/.UYJ@�?�^�1D/�Z�T��]�z�q��M&�ͥ:������㠄�ƫ��J7���6ñ;�&^\9�DӋ�#wd?�����;A^�BMK�Q�[ܲk̐�O��J����F��c	�W	oBw���}y>�'�y��M���	'r��Y�1[�8]��r��'����8^S��������'������Ʒ�z��Լ*�O��X�ѤTH�ώ��&kC�f?ޜ��6�M��>��R��wL<�Qަf��e�r
���&�2�����F	�z�~Ѫ�����'�rB��(�C�ZO�h?��=�P���$�"|��}����C�R�sJA��wq�� �u�Wt9�z��,)K��AW��vN2����n��Ԓ�.q0�ӑ�Dn��:��yĬ ��'�R� F�釢NCՠ�iд����d��D �x�B�Λ����зغ(p�y��Ah��ܩ<�h��|"���z2��x�r�����?T�fkK3i�Z�@�/�Br��u�4�W5�Ӳb��L$��8@�+,=�
��jA����q����;�0�C,��!�ۍqveh/U����q�@<��[U��kL��i�C���9��Q-5˯7����� �Mh��l��&�	��	�퉉�0V�0){yyQ�Vx���h�}��J����'(͈���"�"���!Ʒ��3S
`��9NKǭ[�Ϻ[����{�N��Q�� ����5�[5�덼ȭBqFB�H��8�Nyh��ɉ���g�N~'���W��)�5���S`���|3
��D���"�$�fx8`|�vcL$��%�g���C`�����_����W ���.�[��q�\
m/�\�Ҕ��x���~��GK�j��|1ϰ���1����A�L����3��w���;@�S�T��,������)���(�UQ������ݳ?�*��k�L},�mO����_J�Vw1suu�Z�o9C9��H�e����l]<}����˝�vA�V��IqU�w�,���5^��(������%Y�B 2����cccs,	qc���u6�x-~ ����1)D�!���o�:g5�(I�;?�P���c�>2�$F^�]� ���4t�1��cj�����P�ř�ɞ�3���DJ�/���wuu���qm��B`���Yȓ����ԛAىz.MK�T3�͏5!��b�Ys5hDAN����gXzEG�X�kĝ{���.-��eαh��ȵ�򱠠|�����533���k%��n����W������_a�!Njk��0\[��94��W@ �ˬ�,h�>��RR	����%%�%%��>o��I^J�k�fJJ�2�~`���aV e�#g�ZԳT���$Y��!���g���ܸce����6�=1))�W�u�������F�I�>����}����'�����.j�a��Ul��;lX`�ƥ���V;;���N��n��n�s�ݮ1���1��1�m?p:O�E����O�{�MN����3�4����gS�D�i�(.��)��-!%���.���O4ɚt�n��
o��>=z}��j�S�!Q�3�w���a�IHJ���v�����EW����ʆ�݆� ��]�òRCsA�1���J�'�t@�'�c��론�h<�*�B?�'�P����ik�^0Ė�]77��y��� �F���Nr��x���f���C�&&'��ך}~�����}���i����0e���NjH�Ϯ�L}�[�0c�z��1� w���[S���Jw�z� t��_����x�D(9;;+s�������f`Y�̀dƵC�j93����'y}��I"6�+%�F���{7Ξu���[�#�U�5T�����zc�_��L����NiӪ�f ?��񷂙ԩI��2�!�7
���LD΁�1�u�����5�AW��Ma4k��x�ݷ?K����|!�����x�4d�����ࣥQ��і3��h��\��Ly�]��G�#���L��P��2���"�`�֮�X,B�`���:0�Ź����"��d����κ0�1d栩RD�,_�'��&�p�Gs���˻8��.nt��S���'���Oeq�̚2L�XO�ۀ�8m4!2�p�D�F̘s���b��O�[�W���\��|�<':�xH�u[[��wofM�es778����m`1��T�D�1��Wוo3\w�������]� ��5������V�+S��CzĊݧ���|����^�a���].U��e t�
X^��o�pN���������P�1΍����H߳%J��@q�����+�պ$�9���ۣY+�6�w��Qv^���n2����w�3M��-�[!�^��x�'�����r�� )�����c&�ń+�<{��� X�%S�U����MK�>��
�a�4�o7fO��{��
��b3���CƋP���<�s�=Q]@�Do���j�3���9�
i�~����L�!8R�c�+[^��'K�?���0UGwP�@��u���:�����M�G~n��C�����ɻ������n)Y
4�D����!��b��=<�Bm>�gmgܿ�P��܌�}�@s���$�-�-��X����~�>���z����Q�Y6vv3�f���}�w���Q���-�+���4!���ZZX ��yd���P��-��X��G���t�\������j��+��|-��G��Y���,��\��!�L6�&��Y>� ��7JO��{K�Y.�"��͠���%�����	s׋]�Э���+"Iq����\�=�����0�q! �-�#���t4�zޱ�y��&t�[U�Y%	�d���5O��� �4�/�1�S6���J�i4֭`�����mYF�y��?�rR��^�Y8��kwW�Uͣ2��l�	Qh��'�����3���嚞�4o�d"�t1����h	�fs���4��1��,薩��t~a���u"!-���ߪ�bH��DC5�o.��ŕ��#���=O��7a������Eݧ(�^*0�zֵ��󞜻�/s�H���6���
��~9�O۔��m �2'ɻ?�X�?�i�Ch�6|��Ӄx�����q�`f\ӧ+����bzd��|J���P��-�
�C8Є(
��%����m~.�A�����A'����W�>c"��K���.0%+ ͉�E��l�0���s09qM�O����@�|�SQ|��- �}e<E� �0WԮ�#�0�]�E�V�e�6t� 	��z��44L�泥��is}��Ii��Z���"�g��� ����`�����Xo�� � ���o"�!�ԃX
*��F���Φ͂��3��>�d��_�JJ�}e��'|qhp�;���x
=�p�!���!�QB���+�>~�^�C��B�B���O�_���� ��c��-:�g�"4�w���V�%T�7�4��'�Yx��{�#��y?�v�.5��3C����7751����hH�n���|駉<�޳a�J@@Z�0�ϊ݃:6G�U���?3�d
5<\/�D��?�]Kt�+T6D<��ND]ݿK���***kP�)u��HII�����8*��S�L%-�;���kSt�s��Ņ�{�W;	�o�geB��)[ZZ� ��ˡCw�v�C��k�e{�a������QM��� '�S����s���ixB<!�}��1n�1��p�C��H�b�Ԛ�Uͷ�2@���Y~�3n��tT�M{�[�j�؟?jಅ��5@Z���WcF��S?��B���z�^B�����Zv� ؕw᥵�}*+t]q��-J�L5ef�z�W'�ð�z��&�ե!֊���w���~'�_�B�i��ev^ޙ�a�E۔_�?���c,��߮�JD ���&X�v�fojk������1�PZ���0	--�l.�سQЯ��|?HVGwZcfP�=E���S�2�[�Ɏ����a7����"����,/3��d˗�;\���!�hy�(Za��$[�(���i����C�V�@:��ꨠ���U��we�?��+f���D�����*[ #��Y�����: ���8I�j��:����f"D��`>��ҋ��G�C���G������7�}����>om��g
�l��џ��0�ð�^8z!���e��G9���5C�"�aCp��c�����[�0����0�|��ۋxbz;�?��:�e)d��c�9ݥ��R�.��Gc7�lu�P�_����S���k˵h�*!]F�/J�ʥ��ʹ�9�q�IgS�ɴ��}=��d�΀{ΑwK��py�E�;�.Se��<�2/��K� �Mc$QF���Ir�����M���2|���3a0	ʁ�h\B�d�P6�Mv�w �S�s�
z�D��B�0�/���r����t��:�4���&�Z�ug���S��p=�sߩ��AK�P,�w�_�I(!���/���F�Qk����h#:!Z�	���e�������7%��:���U��'��@<��}����6��&���F%�H�B�G�xȵv�;�Ԣ3�aj+�2��8y7��ҥkY�J=�|�����.���ܹL�!!b6m��hT��<���t9��g1�����rب�ژ���5�b������@x899���ŕ��x�f��K�=�jާL�(�fe4�?���������y/��'�Ѩ�$Mg��V��^�2R\�!K,ФZ��>UHu���LbQ�$y������x'3�(i�
���>���]O�wc0����
�Aq�:N7�w'Į8��#�/��LS%�,�cꂮ4��Ȼ<Z��<�� ��!�/����%A�Ů62kӟ�ԻJܲa�-�d�yr˱*N���V�]���rK�G�($���a���X�)K{���iX�y]vL�O�'�&BJ�Y�t@�Z<��`0�o_
�(�Z�f��a?��W�����U�3�|V=*��Z@���#����!��c�����*��t�O��A��(qs@�LZdR�*�#�F�x��(z,�,�ʣ��o���)�����T�<�k�TӤ��m��ȯ[�f��n�mSދ%�Ĵ�{�gc]�Pļ�)r]Y;f�U�R�����NR�;��Q��"3:ct�N�)��V����}�(���!�Ķ���Z������,,`��W�*�M�Ld0 D�:?�ZDG�G����~�P��"��b<G�i
̟�����m۷�j�we��PF�3o��:s�����+(8�=�'>N$�^����ON�qy��B��$��/��(0��5N����'?J{���9�����-Ӑ����;��� bۯ���Q�Q�Ι�bN�����)=�Ȃ����
��ٯ|�&b����FO����������
�Q���R� ���o�}=i�Bef/wji�EѠ��r&:މ��*��M���0#�O�����9�%,,L	�2�g,"�}�����>���,/����F�)�o'�Y�{}�wO��1_�;7յ	L=iXd+���~+� r��^]p��&�N凴���C�H�{�m��4c��[� �]��{���m�-� ��5Ch ��L<��71>�I�S��: 4q��ڡ�\t?8tZb"O������fMyN
+��B� ��Jâ���!�t=T~���@ZϮ���4>�i0����n˹��3ks0GE�1���;H<]���p�;��=4*���נ��2f�n��2��:��.<G3tī �܏���q[�?��!�8�@<�z^��4�[��PX?'s@�F8�ൺP�3�
�6��󲫫k��6��*���KU�\��.e�6uu�4�Jm��r	ř����@��_�R��I���I ����_�h��a�^;7joΏ�ר��/�q���ɮ�����Wz]x�D}6���v�jm�S��]˼��#ܣ�}P-h��bC���1U8#�7.�"oM����T6\˺�ݢ�t�� NS ���2!x�� %��rY�ܚ΋�IO��7�/�B:�88,J²�R�+@����j�GY�_� �j.e.ۊ�1�Z�u�oLi�!��0�mv��۫����$Ry��B�VMU%�I��|�>x�c&i1on�u|ܴ�jL|�>��Ya����?�kO�hn�K����UofN�H8~<���Ȋ��e�Ʃ�eܐ�sn�� �}M�j#�7��eo�ذ�%��6E���ㇵ�e:x�2�r���E�[ˉ��\��v6����kn��w3nk�Vc*
Ŝ��y��u�Y�.�q/f�Hq�7L�0�*`ב<�W��!kh��K��ۈ��;��������}7��K��,��e��i��ǟ8��f��y0�~��;w��0���7��'My|4R-=1�3�H���x�P��̙��ې]�[G�k��l��q�~91��w�bu�����7�����0��~ҹ[�1g4b$��Bi��l��+�+}��;��걅Ϗ�z�l+����:N�ARnyKߺ�Õ��w�
��"�\\�!���#S���Imy��b�T��N?6*�=T�0��B�BȌ�|�X�D_q��|*11Qqܥ�e�@���(�����;�\��5ݷܮv�1/2�&�����0X���	}������z� Ϡ�נt��a`���;W�O�q�w@�f�=`�V0�L&�a�����_�v�z$e#ct�EiVE��Wsd�e�gN����?�߆E����Ӡ��B��#���o�>�m9���4�3�����L2ݩ��#�.��}������9E�6�飵@�(	��6{�q�����=�Ոәak��M�մpJ|�!O	�j�G�[���"5�m��zĊ�ʿ
.��|oV���:���N��;��#���c>�~��\Vw����K̗m�S۾%:�S�Y�ߡ����p���0e��;,� ���������|�K&��}�/*A��ѹe�7�gg�G�Ummm�wu͇�~8XdȎ�C4�"v����S�4|7�A���5Ο�_��P�0�c��󝪥��ê7�r\%�w�IS��}�Y��	)?�*�a�qe��i������&�q�C�t���M�*��v���@.Qh---����r�H�ǭ����v�ީ��Ӯ%#z�.��<���������Qf}}�L��W�4��kVV���¦}��s�������t��IMM�ɪ�zԻ���ݼ~������S5�S�x���&��uB�`�B�q����k��~�PO��Ib��Z�x���okK����Xp����)�5������1oR������F��
{�]'�N�,z������a���	xò���",��n�x�˭������p�T��i��Q�V��#�n{W��T��@<��Y��&�T�?�h�h(}���݂�J��i�$//ozvv;���{x�b���5�����hD4��NM�^K��_i+linN���uȃ����Q%1d�⌃��]j{���7^@;K�����!;rv�*��V��t
$;sn���ׄ�������ޒv�X8�zܧ<r���u���_�/�vq�￷��M�L����Ӓǣ�~�Gf�fX����HOM��ļ&����~��)ZџT�$ZܡMz�4QW�Bj��Y�H����I�1��*ʼ+�lڄz=FcoTxˎ�ޛ]��y	B��/_�dk�����cQ�UU}2l�{nap��6b�x��P�d��� P��8O��F�|lQ�*a[^�.��e���g����~�`}==ކ\�u]\g�ōS?�vµ�������	뫋��Z����|�:��. ,,Ɖ
��AdN��\<T��{V��]��&�`{��lqjJ���axܚ�b"{w����>|�9�+?/t�p�~zz���0ͨ��;���'XJ���xG��lQNԮk۱uK�Y��®�i:)D֊%?�yv]����R2��vNb!�,t����4��:VOBn�Ϧ����͌�ӴuY��� KJB�X]������/S���pK��0�AոC1�|ӄe��LV���%��c􍂢��=|���!��� Ъ5]�J=���v遾�G���U��.C#�����Xk��|ic�'��?���B�k��D������PK���{�/����ٕ��=a_�]TQ�4��vڌ�}�2>�Aj��1������1��>����/�{��OX~���Q�>�17���:ޑc�lVIӃ�t��ӽ~}��l�s0�lt��y6 ����(��7�	����=��a�ǩ�$HBԒ�4������=hE���C��Rz�	��VVi�6Zx�pp�Ȑ�7=n��. ���&�����*Nl�:t�i~��N]��c��I#(q��b_I/ƱZ.�z�֘�'Pc��<�®��VɎ�����>���N��/��Ao'��7��E�d3�h08���lvf�wgt�JhzFF��n��\��q��.�}���� ő7ml24�d���s���g�Yx��E +�W�&���e����؞��t���Xj?����yLst��,�>7�q�d�E���,c$C�JJK{rl,������eP�ӳ�� �p�����b$�I/v�J9�N2F�P)�ܭ2�K���u���<�Iː�~��p�9ckc���N��\[��m����������kT��{���o�}r�HC����W���ӸwZ�:�w�Ľu�)���~���-l���~YLL,�(���qr��!��i�D�C:Q�?AN�����o�f�� �UB�ij�Bb�-�T�̑
< |�ON�:�n�$|m?�J}�'��믮'J�8�����!��S��.֓g9i���gH$R$:GIy;yq1#-�+�1��F�I���ߍGϝ=��!#8�_rY�61�3>�����"0��]3(�����s��s�8R��I�^I��ʭ��\Pĝ:j��eBŨ�aNw��8�����Y6�?+�//'}4�c �~�	dmE����'��2q�c����d+���J�4�/茟~S����v�{���[��ye�۬����u��V73!���	��7��(���J ����bN�>�Ȍ�gd]�g��gŰ�^O*��S��G���Ԇ�%�(�]��]0ԑ������E� �1��@#i�� ц<y	��U:{���7p_�'�^����U6;;�F	��a����B ��v%��ϘS�n5
Ī��!�ODs���ƒٽ��l���~n:	�t1�	 2�c$�s&�ϝ�b�3��VT�]������-A9���"`h��?�o�d_Ԫ���N#�Iu
>�46G�w��Ԏ����А)I~�
r��}�vc\f����W���]0�&�9k�}o�܎|4�@����D���%�y�X����'
�6,v9�?}�{�;#�zΧ�	.�{B��u�:�V"�&�+���~	�P̡O�.�+���Ǐp��UB����j%��R=JW�hS:�(-)-O�~�lmcsĔ@��hG�7��F�9�6j��_^:�a�yh��ڒ20*��{�:�^@Ù�\�M)+3�v#���)�ʵ���b����]ب���L5d��Ɔ`��sM�x��X��#�y2�7���K?��d���f��wt�']��A�7��#{�Z4p�ʷ}��h�oK�7�jsD�z5�4���V �2-�w��MMb0��;_Tiw�放�k�'�h ��^��8�Zv�^��k���K?6��ʿS��+B�NN9�+yU4�#Yvl�a�r�nn� ~���yŭScKꈕ<NV�L@=��v�{tks�0�S�_Z��UM�]�n��x����%��t�x�;��,v>�����g��IJ.%���2�ί��^�*[�a�P���[j�ݺ 1�|#�~�xTt4�B0��!�7P���T;S��K���i�s	�Z]���X�<�Ǟ�G���6�}~�w/���kIj�t.B�iR���QN	�J�����0A[�?q��.��*%�J�6{��+�I@�ED�&]\>�ά�]�^:�x�lz�����J�m�Q�n=�et��{���]z]��RS�@̶o����p��Ŕ�V�a�J��V>�&�	M����%)F�6p7�	_�mw[�]7����%�h�/����F�ݤ�	۾R��!�f��b�)*>D�"��&^��}v��`H�ܤ�O����<�d*���w��������ovu�*�L�:�Ip�s�31#�����������e7����>f�Kɔ��k0ˇdX���/I�_Kv���P��2ً��f�8�tvwgTl�O���� ��۹6��G�ШI@.�C_a��w��ml�([!f��**L���!}Ͽ�
�E���Z��{�&���С8!�	_8�e��QT��$����/�"Ta����&��U�/��'/���w����v��Mk�~	*k|t�(�(�c�iR!�Q�c�]�J҇����J&8�������Ŷ�:���q�Q����~{�Y](��*�4h��;�]<#!�ӌkBS���L���V0�B<o#�\�uܻ�@������	z�s��rJ3�ܪ�����|������d�����)�������7�-2�M~a�D�Ϻ�Ŷ�?˽VϞ=k矵�:���y+�W��cv��c������ַn�P?�p廽�h��/�?��:Y<es֡�4�}>n�ޮ��QI�U�JZ�/��/�����F�l��Q>&�a�����	Mw.�E�022���BH?��2�aia!�~�,���tUP٨7 ����`�{��⒒֞[�;���Q Q(�F�E�V�{!%-�o�+E���X�s�#$�N���9)����S��z]4ح�k����;�ۧ�U�*�o �wǘt�r��A�aT�p�0(�.0r��6*/�v��{ Sh]�M�Iȋg�z��8��,9X�J�qrr����$N�5�:�s�U�I�}����`!���u*�����L��Q�T_�a�u 7��\!��+��旴����޶-{��	��3���yu:��N��ďX�5�q�G���O~��=�g��<���+���+�S��Ǐ[R[8�BY�8��5�^�Yt����9d(���9e��A�9Bb8�������0���﹯㹹���N5�t�m�0c��m5�3AY���+R���ٕ�'t\��#)���:��ل�{Ĵ���?~hն�jMNNJ9=B�.�I�t��6�t|
�K��KW��	�JG������AY��F�b{�k�l�F!��50HC_�K����6i�40p�b�,��q�0����,�X�C��^n3A1p�3�$����kU����ME�2�8��TA����h���V��%�ƴ+��k_��AF��M|Rqp{�@V	��μ3��&&�Ku����b�6���A�bCoUmɄ~E�����yyy��� �kmk�hr�h�d17��<�\[���r:��m<!��0N����	�����G ���|���׭�8є*'А��B��H_�����C&nw�\Ҕ%�3p������9�<���LK�>�������ҋp����=�����I���U�D۶3�M-N��q�D��$��q�1Eߣ��vB��U�lY�.���|����@h��Y�Y^����d�v�!�r�T���ٳc�)�cV�Q^P���J�S\���x�h]t萉�������gr�l�AWz�k�zD�N*P�m�`����/Q�FS�&ｆG���*�ӆd����<w}&	���9�����غ�6S���kn����vY@}�ÇǊ?��U��s��ќ��/��v������4�`� %nT��]6ْ��j�Lsb��vϳ$��ʘRwN}��칟�/B8����In��J�m=v� 4#�'�H�b����@����<�Q��~'����m�����}=�$�u��[�)Wߌ���u뷳]��f}&ԧş˛����H�a3��#7�o�t�_��4�@Լ�&io�T�	!���7+��77w�NzO�߳{�Z���lo������!�.g`�6ȍb��2�0��iEYr�pwg�X���+*�s&x�.�}�1���w��T�@��24�x�ik�ݖ�=/�9'/�4��f��y������������~�u�2���.��Z�!��`�l�7!Jb��QܶE�&^+Tf6@��4����:�T4:?� b�4_^.����ӯ����/�2�.���ɫ@�+6&*��S�謔���͠1�>"]����8(3]I{#��	t��%�u�dED~���j����E}�`�`�
�2��phFV����������N�Ǐ���"cǎ��C�^�ꖖ��GR�m�鷉J"����̻�=���֤�{��Յ�kI�v��,����.������J�~����)�l{o ����������ב&;r�v���If-}5��]�Q������N�̿��2����3G���y�6m����^��(���)�r	]�
��NS-[���}e�.���8Hb`!�<?HR�t���r{6�?<4�g��xcTr���wf}5Y� ��Ѧ=k��j����E���Sz0��ӿ�
�Z����7��K�>�Z!��(�?;����Ϛ;�yYH$�A�>R��&��x��FB����;�j@� ���,v��'D�6�����\Fcݨd��(X��������^����nvβ����~��z�x�gتfh4$a���NJ�q��� �����B�Kxv@�)��py�`���.���A���#����թ��B�}�=�����$�5-Lv��4[�X4=U��i�HM����֬�ԁ��l.8l�?L]<����R���U�d�SFI�(Y�d��NC��d�B�=�*���/�${���_�������o����}�������<���}��C��A�}ʀ��9;?��%�|P�m++�v�!�B�Ԥl�S����(̾��0����e�W���B�Q]CG'
L�m7|����1+#(�̫����'5�e�n/�^!�;ͱi�cz�j�컌��c�S��
>7�NW�\ǿ��������+���LH�٣�T�>2�d���ɓ����AMM��'l�"Y���sw�%A���'��K�� �׆�����z��FGL,$��'Z9І 0�^D��I�7ekb^<�1a!ہ�yz&� 9/�6������2�bl�V��z�ӱ���4�]A�녙ԗ��YMj��;l���ok��O_�;;�ޥj�Rt�kg�o���]MMMu���|o�����	�6��@�!�����������ޜ�0���/g�}�XםK�g�ٍ����ˠ�����UC�έ��g#�z<���,����>�<�*���3����\����s�
�|��k|t��[�j�../�{�c�1@YȇH�6[9EE"��\]]׆�3�朠�r��`ػ��lmb"D���u�A���-�S� 
l�Q����ZG���o�&C���ko111�>�<<<�V���x�":ᾶ��h��a����KDiUL��;${�f���R�1i��C�l>;T����)�I�m6:�*-}��E�߿T7��R9?��n�������g׮]|g��ZZf*_���0Į���r�DZ7�҇n!ʾ�g�ӆe y�)}P0	(�T/)���������n@�R�F���W����6G�6G���}F2�vv���)] p`΅s�R<���VϋS��m��������2UPx8�E\����o��@^�O���q���s��ԁc%��"(d���	��h�"#�K������?�CA��~|)�Go��$$$@k��{X��f�l�n/o���s�˧�@c ^Whi�Zv�g�zUgb��$R�Ӑ��[e� v��y�����.�z���H�m�=��ϟo[$����)��ю2�\�69�gZ��V��<y��&4��q�Nmm�W���paa!8��~,�5�^�ք�[����΋?L�3߿�ta48�>xX~U�d����zƾ:��(ʧ�F����r;}���w`�gbT�Vf�V��:zzѠIC����ߺ�|n~^��ؘյ	��5=��3HKKS�^m��3��6��bZ�_��&�KP���~;+���R��P�����+�~+��Vm)
�9E�Tvq'y Mm5���TTQ�O�f>�B�URrJ +'��=m���X�G�H�-#��4��YF�3�t��
/��:���Jࣴ�~Z�1�������<�&������D	i�(�Td���@�7=�w�P�A����ڄ���C�f���x�}v�/Au|c�Н�W��"'d������FAjw�d���˽�U3WG��Ӣ�4т*���믧}F$�v#��c�������B�����Ļ ssf@£S(�Z��&^l�Ȫ��)�ܑ���'������[v���H��;�M�B�<�ୟ?vvv�zƭ��x֣���@<ȷ��`��7�ݱ\��ak��M8�=2.l�����+rE���_��U��q��뼼V�g28Fz�ۥ�� ~�:����E�qq�$_--�A9��-���q�:��E�v��-@@f_S�k7�/�G�Qq�<c���ۄ	7�H�ŋKx{�/��_= mo[<
���xT�Y�7㖦	y�U�:8D��.���4ӡCV@bE�9$(�B=�rE�=.MW����[�#�A���Q�O�sf�5@#�W��Ց�U�,_
޻�j���������������0��y�zy@y�t5���޻M�CeƄ����2�Ъ�/�ƻG׌�����#N��+�����D�w��B�xk�t���ih@}IK䵿�	�ݒ �g	��K���Sﾟ~��f��4͟oo�G����ܿ�6����ꆆ	����iM��%/W��ߖ�nA��!�clu��w$/M�e�}¼�p��{WE���U��e������B��?�t����Q!f)��"��H��T����־o�|����ȕYT�k��Mp��G�0�"��OO��ȫ�D����`�(�4ʥ�<ڲ���� kNN�̩О �{��H�cP��h�6��,au�G+��� 6�ٳ��q:ٺh�(�.Հ2ZT�a '!!!��� 4*P�w7�W� �Ҕ5!| �hـmY�~�2�,:���֭��b{���F�@�뭷�g6��u����^F�IHd�o����iB�V���(k��h�DБ�'�6�n|�۸�� �{U<?�Kw���pEة������{z2�d��A�A�;����zun�l�wtFs	Z,�ԡ`K��N��G�����;�w�=-r3��*�Z�s/��N�z/��g��qR���)��7;�� �>$�ms��kt����2�j�>�N]���Uѝ�!��^BB��8zz :`h�vs�����E2w݋����
���룖�:H�v�
��oLN����@�����G
]�u]��bÈ{]��m�:�%�];.;�ٌP�����wZGS3eu~���x3�����]�k��~4��ٕ]����`�`��S4k����[2ڮ��r�W���m���Toi:�)������Z��]ݱ ��o��_U����T[��ޗ�֟a�w{���*��r��A��(�7�߳ �}�����|���?^K{/��Ӗ*�܀6%`T��������ʈ�f�����ծ?��YJG���2�1�#�w&:6:��_V����¦�g��������m�Z?��u����x?�+�ohPd��P���K?.����8?�J^�Q5<2��l$�,����8؍��1R[�����@Pi������۷sRh]�f���
��o�AJJJ��kPO 6�{O��WTH]K�1t���8
�
�����Q�>��ӹ�"^�K���n::��,p���'�^�6ݟ�NM�qH�������#'v��0${�ƨ G�ƭ�-� w�ϟY�ݏ�"|E�ӳtllL[O/����
�{N �k�S���mF��;8��}�f�xn��P
�&��,ޣ�"3��ǁa�A�0+PK���U�/�<t�8��݋�J9�@���)�<<���q	?̆'������f�?y�$:���-�B�ڵ���MQJ�� $���\C`�&���҃�[g��E;�g��)J~��������ľ��oPg_[��t��ݒ�ŗ�������`^�II~�ph����|:���,��Lհs���WS7��诈��W�����w̜r����DhiQ-|���<+kk-g�w�Ьҳ���.��!�`t��"y�В���Z��wEЃ�����+��X@A9�5��@��Xm��ZxH��^�SC�*����ɑ�̣��KZ2sz���%,&&���d���jCR.m@-QM/\���:Qٱ�� ��I��E %h�(=4 �+���:��|RB���N���9���yM��))ǚ����l�{�Jsf�ff$R�{9����EЫ�M��rؿ������w��׺jj�i�AZ��|�HTd�t雀�@vff^A'D ���s��ǅ�¢O����sss`n�ϓF����-m�a
��|���$yYx�ẞ�kTn՚UC3ڹہN>�M�EE���I|�y�ݸ�c���%7�l��ŝ]���P�10 6 N���!5ŧ�_�[_����K�(��F��l$��-��A����M?ߵ�+K�'�x(\�^� �"��8mW����0D.�3T�2Ai�=��y�a	aE�
3�z���p9�t��������c�ck)ӓ�]G�+^>}ʀ���%np	�t\)��ȸK�{����W��n^G� ���'�Q�?�c�����3�`"@����x���?�t�+l�.c��I��Q�o:6��oXlH,N�JC�����W�@[��������2.��}��
��x���6M3�Ï��)� �c�I*�KЯ"�T���nl��?��l��}DԮ\�6��'vb�	:���J -{;4��`6�Ç�9m�4(Am��(�����P�Qʆ��@M�Uo�1���;x�p�X���ΥK��w`�-d��#���.�j:������<�}n�IZ[���?�V***f��&�I�_�H�KX�FGX��nO���������2\f�2�d�gƕ4M�ʧ�eO=����售)х!�No3��F��=9�����-/��t�V��ֺs�K�5t �쿰Tdލ���H�*H��Ck8��oK?�?�M�DI"A��1SV+
�=;��: �+��@��h���j�lęz����t���wٰ��X��1b�[�����x������&��(%�ګh�z��3��w�&���|$��Cx�b����������'�����((>�r���о����<������4fcP��VQ�S�S;xʝ0L}$b�����3����R���i��/���Ǟ<~%����>v�T�,������JF�.��|rm������Oķ���B{H�IP|���6��M���_��rF��g��+���_`Շ1OT3P;��:cT�j�V�w�,�C	7����;�3������F�f4/��h/((������>Y�����ش&$���^��F�N��`H\��e�#����.]�Ip����' z��)���ȗ]��m~~~�ÒS��C[�))]N@�]De-U[dk���_�n�C���G�e��qq�$\�	�Rx�����{B���u��YU�/@��E�^�Uݚt��<.��"6?�aZ ��LMo7��;�-������വϲw�W5p���w��*����ځ�.q#�� �\�^���+����?+�PǅO��%L�3��QSG&%���K�r�:s&�}%ZAE�6��x��d�[����V�OTN����z���P�����$ٯ7
��NJ�,&!�k�M����īfT�ch,8=�E��g�c��F��^�>�2ɟv|6C��9|��S�4'a�������)��?���8�D.���ee	d��%�R�� b�*C�zݒz��	� �T�	�%mXl�oo�K�T�e��"7E=�D�SQ�i�*�xG�����`F����3c�����������P��X��o���46YL��CS�]>z⿕G���is�>M_�<��12JQ�|���O�z���N��F�c^�?k�_ZϨ�6�"ڵkW"?�����eb�8��W�\�e����V��ɟ��N�.�'��o�׮��,��������$�}0�y��Q�̯��u��隙4���	���9_u�������+o����,��35�M<}Yh=Y�D�/JS�p0p�Eύ��������u�h��ߛ�ƫ�@���		�����"����;��E{����EԒ=F�]e�;O��͸Q�'���Ǐ���z"�L4���1���5�����0'�٢%a�v���L�-�����O�R�e4�B����
�L��Ӷ�ݐj2�um���IMM=�ʪ!|X�4sl~%�W�:����ˉ���u&f�k�����Kqp
�&@�KI��<8��[�A��(>�d��ߴ��Ձ��v"@�`ra�g���� �Z[��鱔�6�ܲ��\���F��魹�y&ꇌ4���jywz��|�Qy�;4,,l:(�<0`���_�����"�ز�b��2z7��}*�nC�Lt�9�8r�����Z���x���%.�2� u��6(���=h��Ά��
3KRj9��>V�^M�C#:T6���ڏGI7���9��b�[	p�@Q�\����htad��itw0����I[]ݡ�V�^��%��-�`@�p5@�~;���ˆN{������E��A���7�̈́�8�b�tμ��0 ��7X8�Ŝ��*7yR	�5��X_?��C*��p�]�&ڕ��K~�.;��F��K `h�
iS�yr|��O�����U�F����#c��+�X�)�����-Qr�4�����
Y��J`��,�ٗ�\N_1�p#Tz���*U���J?y~�L�N!�����d�~L��:���r�����}r����P�C���������Q��bo�&������*�v�W`�@��)�^����~^��v4@����&��[��t��ꀟ���F���"F%6l� +�\ �����	�oѦ)b��~�v��r���=U����F��AG�B�&L��D$]��_��LC-B�>��|f������;�����_��=%~�f�����;�a�d��|���?�����o�ܻ�����6�dA?���O?��X�@�V��Z��;�������߶x�mll�K��2K34��P�"A����ߎ�8�D�3m�!`-Z-M��w��a�)�.�ultT�뀺���}�B�G'&�+�:ٺhM��	�J��	�MK�$oTAH눩6�=��1�#woz�*���^VU�짥�z����l`�U��wZ�3%�+��qP`5�^��������m��3���0�:�H����&=���I�zs��U���lo��DOE�탎�Tɠ��QQ8!�C'�"�6BR����l/�>����ӧ=�V����́6<�9hXtU����h���j\�� �&+�E��͢mB�<%�2I�	�����Ю��@��?�!�6�r�࿃����d�o��,�^�M���/D]ġ���2�*5Oc^p��I���
�&����>����]ǴAL򒻷?����/:_�N�'z��BN����@>�xo���;��[9M3=u`Ghh�-�;D0�vA,.�Hy��e�g�g�j�Y#���i�Y��ʥ��g�`�f������C��QǞ�',�	%���0��ˣ���ZJ�fs:�v]�u�/����!�h�}��6�f;��<NÄC&�,�6&��
p�7@\k_���p����^;�H��^zr���xH��$%%��� �S���P�W��D�MO�����"q�o�RE���]�t�TP�4�s$B9��@�kii	�f?\����WXo�aX	�qs�nG�g�;���J��sfՇqB.,���G7�6t�A�9���ȱ��_QϟKl�� ���"�7j̺9��O�n��qVЁ�P����|�V�7�uD�ȈC�6���گ}�旒��Pocc���������eۻV�l�hc7xm���<�9��q�s�Ɋ�ᐩ�)�O
��%1ee:��<h���>0���.�8�m��y`�n.� F��X�}��/A\C;F����ol��ژ��̒��hA&7��!�9�}���G�:���V>dA�-��kql��l%�C7�t��g���|�I�A�C����mmm���b	�x��v�A�ƍ��������--��9�JK��"2��S��Q����ת�Ckr��ţ����"y�j�x�w�	����ǡ|�r:�r
<*�L�E~A�I��[r����	,�m�"�q�B�ܹJi�\�}��b�3g΄p����-f���.=cs��ן�Lj�NjUZ��u�!xyh�vղ��>�--�@;$
��t6�D�u�9���T��C���qn���!����*�<
���	� ���ח��o��٫����k<go���� ��E%�dq|N�߯�د:)���4�Εhh���N͂ꨭ�3��̼�֑$��PP0w� �<�>���qaO�}d���d�az�;w�
f#̆m��v���	�V���`���X��Bkv�E (��ٓ�);�-��,,��'3B�&'�R����=}Z��Qgh����LXPPpP-$�=�k�.po����p\��E^�;}�<�I�U�K���3��Q���D��$;�D���x@�)�������F��Q�C��^��;���@�$1C�� Y��L{v�4:��_�!�H�.�����Z:� ������[]����P_\B��n*�0��fu|������+ۿ��\�
�R?�xЩ�-�(~m��ML���?��p���oFN���k�����L-]݆�-�ĝ}}҃��¢��QzF���A����LW`{S�r�)4l���T)��Nno#����Qㅔ������EE"(g=|>�<��X[��-�����7��15V�4�j�"�L�[G>�h���#���jo�$:�x����q�IX�x��l�hee%z�;X�jJD(3��E	����1�������	���v�mmBG�A�|�<K��DsRTRk�~���9��� iYZ��O�|v���5чw�9�9�N9�$ѓ�Y%�J���Bw��ff�����ʇ{f{T'�0~q��\`s�"�Q��ν�-;Ξ��p�sfr������}W���@������s�U�����|�F3(/Sa4h}��fq��X:����LB�d�U��.���8_����5�E�_��
;� "*���͕��5�|X�2ڎ=��̵J(k�;+��Oc��I(/UU�(��ΘU���<�<::�(/#�Ay_iyZ�]�Ԃ��W��p��P�r��sX�Jh'T����P��|�(�۞#�7<A<A9n�(^�����\76���Q��H�@����ﺁ�T�J5!|kyk�xbj�Av�(K+x���Ga"�1H�^D���(����	�{��1C-)���ϝ�O�==�`��s�jNtD���4�~3�&ucG�����ꍜ�Jy�Զ�2���={渶0zz���O��#���������<fo��ZQ^ޅ�Ă���bd>kp���u�~��-�Qޠc�B_v3�}��n��)EΜ��fS��L�}/�=��4�ҳ6�-��v���r�i�����c���}�=Y���&���?�:�=S���~�f�O
�ډ	��N-���!䚕F�\�w��ʘd�V[S����b, �,#-	��zy�aONjMb�Fy���q�Fm5~k�C���P�.��t#M����=�,�&O
u�
��caA�s>*�Ϳ�vz�����skAm��fA>� y���IU�Q#��Z!e�=�r��e�b|hWW�]�8*�p�+�-�?�˱�fL�b�� �;����xz<����x0�{�SZZZ��':��M}}�9d|X6�����a�h�0�8�W�ij֘놛�.]�������e�ǭ�������f�֚��;v�� /F�C6�9N�n"�נ�T�/�|�7��ҕ;��h���p��`m�[�ڼ`IygѪ��\�{�$����Q�9��<��y���ahss3�auY�a�(H yt�S�)h/�'���f�xcrSA)�M����m�g9r$���/�r���}�,*�[AZ��of#��2@�:�
fJ��ɹ���5j�I3�?��FJ|Q�c�}�?�s���Q&l�|�^m��+����nt�"����Y��m1>���!Au$0��yDU
�9�jV�����3m�%Z #���F��l�l�y߾}�c��M��F]n���d������~1~F{�@�;���H}�P����p�O��|]g�6r3��yh�VV�y�mR��28Hvs6|��{:F���{H�kew��5zWU��!�54�kP�`_1��7���0AN���֗�����NtY�>uF�����C4[��@
��8��Uo�wVx��.�=դ�s��0��7�< >W^F�9	�aj���$Z��vtt��۬
o��^��?h�L"l�Ȭ�G�_�|�GQ�Kr��tW���N��S�`l��h�t��2ä����n
~r�`
�z���)J�լ�>��-�¢5�w��MC(��75�)���b�C�'e�$T{��e���ky���n���F��a�iA屵74(���h*��,�?V��B��wsQM�a���L�1���L�ꓪ�	Ӎy~���o��b���i��, �����>��V��y���l0*��U�r�^&Aq����u��f���C�Z�,ۅ���g� ;����XQ%���x�qFOݼy�T%��E��=E#�A��\\\�j��`l�+9�EN�-�Q����Z��Ƹ��699�"�5�%���9G�0�[ZI<�b����{<�SrvvF���+����I9z.�d�qw�w`�K� q�+;�4䤹$�{�ڵzT]0G�w=!t�S�EQ���@�<������|6Cv��5$_;�;j;���M0����h�fko����i÷r�=��l9a#��6��Ot�6��mLX���?�U��L�rMA�nn����ӯ�ι�_մ˶�>��,A�����Z�39�6@����P��bT��z�*���L�l��?�}�A��3�<	�)��܄:���L����/.��h�.�C[#v�����U������	i� ��C��wމ���7n�&m�k5���*�2��Q�pl�����R_������P�<�U�N��If�7�3��x�ʊO5A�)T�k�K+2��uv>ߒ(-�@���δ$�r��Ae�鴺 ��Z߾}��v��@���͝�v����S�����o��
� v�Er�U���U�~�����~�K�L.lt{�{��?,�Y��3�S�������Pw��b��j�We���(�D)V�+�U���YuY��s��<2�H���&�E"�csu$?�vNJ ��n�F[��q}e<}�����Ͳe��
��d����Ϙ�O/��U�_����nj#|x?L��/�����o;:
m���/�aWL�uO�c��!'������{%I4\�	:$n�dT
�MKK�z��j�FZ[�Xh�zIy��N�w\����X���S���M+7釲0��Tkkk��_/�}�����KV\�7h����l�+})<6T���Z�%F�������N��INW�`{�H���Nn��n-%�
�����d'����{@Xk=(�1��ӳf����#ܪ�G���9;�K�g��P�߲��(�����0+�Rd�)j
u���ń��5!��/b&��ׯ@�K�Zs�A�"�ݹs
2A'�}�-U�@����׈���Jԗ��R]<G����ʏ��$6����ΧW����?���^�Dz�S)�k�Da��jW)���Dh�_��: ^)g��V����m���r���$m爞��ݏ�H����+����Hh)��e���=��� e�ݐ��w��o���f.�Ȩ2����C�S���ǺJ<f�hQ����em͏�E���PLE9R�蹑Q��h���VO������Gaڏ`N�+� ��M�]����U���(GMAG�
�Zl��4����.C�5H+�d��_���/���-"����4ײ��ZH9w�Y&IbQ�T\�I���>mJ ��fX2�@X�D�7�f������P�=F�� ����o�O��껞�S$ b����G���ś��y�K	iRX�$�T��>h��0���6yMv7�˖PQal�Oa�799����72:��ъ�`�0�i:ގ��;�ust� ��%�N���	�^8����&���t��Q<5������Г��$~��"m�4
��q�q��}�g�&��pWSx��1 �l��O�
رvP��b��x� b����;�yֺ�R:Fię�ȫ0����pԏ�^v�]㋯�|(唷[���
�F<�J#���U�Po��%՝��\�~9���hcU��I��(_i��[M��H�ݜ�c�����	P+� 4�H%��W��k��!�Rx����0bJ��:��������3���sr)� ��x��g�h	�9ϴt�}��.�����+���x��fy{{�?���"a4�Dw��Y�x�L�/,����I���������I}U�����ށ� JW�;0��(=����,k�Ù �I���̀��Xx��ܪq$���Ϳ��`�,�������!�L*N�=���k0�r	�"=hc�'����5 /,79}4z���<�ʗ������"6V���79��qs}u'�� �sHZee��U�Fq��9����5�_ �U~�p|ыPֺ�^M2���ݏ����о�Q���S���P�&�{�u0l� �����CFo��Dl��%d�B-���ŋ���p@F`o����&�i��om����(�<f��uP���q>��(e�J �#I��7Uo,�*3@��?�B[s]�}�`��4ٞRc����67��i��㠳�M/W�ͫf��I��*���(q�5(w;nL��`�#���
����\Xl�t5����;1�T*�� ��g�Y�6��6���������P���|�( 47ܤ֢%���n4Pf5��a��S�|����G�ͫ2o��߫��<����RRb[�O�	RV)����@,bf��FY89ҝk|��٧�&�I�}*^��m�۬L���E�9?~�\kj]ۨ�u���v�>��\�ؔ�����R�ŋ��.��/G%���֣�'0h!ԓ��bf��+�]gJ,I�柎󳘍�=]	P�IQ�<�	�x��ԣ���a�e��h����.�vW��?~�4����U�|�i����)Zp��C�nv�$%���@&�e999 &�W{$݇�D�M�䛌�FOR�mƑ	V��G����x���������q�a���~��T9�%O �Ъ �&Q4،-�*����n��R!$]V��yՉ�`>�Q,�ЍP�,\$�Gh5b�����3gP�A� N���zְl��}��E����O@>��։_29@�P�����Fg:��t�(�͸&��`a]��>"j��H*ʦ�cI�����W�-�kX��G	�u���LƇ�n�@�T�H"I���Ą�m�W�Q�y�c>	�����`�j�|m�&����1����E��;�X��HvȐi�6�H3�~On�z^��$J���ק'/bb���jC�^�JJ���qsw?xr���Rt8��$0��L
/!"�����$�� V��=mI&�V��}� h�kc/M�'�N!�+����zv�m�����ؘ���z>�U~:e�(�aL� ����h��b&䔍����ֆ�,�U1��E�V|�="G���n��H+��L�Ȭ?��MM��0>��r��*�AZu
=���"����j�T�ZBi\��z�!�"yLj�2��+[�����J� X�OO����� ����KKY����`�1>�S����t��Ą����k�������Ж�r9A�{��#M���H����
��1�V�Q�Ӹ���(k6���E��H�0��|jk���]�i��#pb��T�Y��dw%$$ln���3a��]ը��d٦�	]	��.yi�M���`J�r([ �)�/$�P�ĺ��o/��f�a8��r�R�tCL:xkk�C���� np����[�l�c�YAo�R`����A>����-����?���r������\70��U�՘3�kcmP��=8��_t5�sM�m㋚���x�:�1,E7�>ߴQs{� W��y��R
����m#B|�*s��x& ��� ݆����% ϟ��|���Z<<��2tf��cRA����0�Eie�r L��P���/v�ХY����G�+�<L�xo��@�0��D�h��ӧTw�MA`#�����ЙB
�/��U�S�7���)�H~�k㖔�g0,��Ǐ��Y����0yŤ@)��U��'Z���`��aZ��������,���T�g�de��L8�J��+ �{�a���|;�ρl���<����K?G���|�h�c�S�~,� U?-�4�ՈevYmsc�E���o���,)�� S�p~<&>������Pw$���+w�h�#iI��p�^>����S �B�}·�k��I�	3��G8Q{	]8l���f*Ŕ�e����k�C`Hz�b{��u�اP �{^����}���d��EOa !�<ת�����&��(�g��y1uv�dڮh	L���|]�ѪT����`�� 	�\���[���N�R�l�ĝN�%qt�� @h�����g�	a�`���+� ���Pˊ��?6��V� F��~[��&�M���I�cknn���Ԇ�[�ĵM���o(������b ������
4@���A��g�F���3��{`�%�#311�*���\ZZZ��$Eˢ�b�P�E�e��������A)�`��4�֞�y�\-W�w�؀��E�KU
����W&&�$|8�ER�pxFo\�����L"�G�][h�(����g�W0\��ʹ�چ߶���u��;$8�4j]]]�h�'����;���[���,4��Ra�<(t���? �=�T�`p�{�0����I,��6��i��@9Z��Z����+7��//G�5U6�j��C��HP���6�n�~�{H�O/s�Bxs��١�N�G�<A6t�(���IN Ԏ��i���-��H�?G���o��`�_[[�Rۀ�1Bw���O��I�R�� z����n7 �,��v���	�ʈ5D@x�
��k`4� %��q���6���}@O�8��U1�j5J(g��=G�,���ZM
l�p��WRqH`�
�9�
�z�&�!���%�R�ǰEk*A�
)��0��i�M��r��JYoFoqQH����Ԙ��}��Jg��%���I�D'B__( ��|�V<��`� R��1<g$Y���A����~�����rw4�0]�̡[�����҇*Hp"�$�����B�B�4�k5�&1�������Ps���
ώ�Ll"�5�8��;�V��$�ӱ�N(�)t�j�I���E:���,X�n(ٻw�mlI����HZ��z��Z��gSe�M���͛Wa;jCPf���So;8�Q�w�o���@���#�9?Қ�ߵ���GY<)k(ؑ7��5��c3��I�Ɗ.j*��a�,���=��:B{i�	E^T��h���4�(LX2a+�d�d^�4��T�Q�&��#J/"�	�x������x��g�6�Z��FAY���Q��jt5z/6�7����<4���}��?. ۆ�W��W7���\f���v�<4���b ���(j7�w��.Y��|��<*���7i��/h�۾����`V;�b�sJ�wٞSc��2y�N�&��F�;��Ǻ��|�y���+��W��L��j��՝�,�J��EP Q����Usu�J��Fݬ�C.3L��DN�B�����;wRж�F�E rn��؍W����]��$3*����1L�� H����"""��@�
#�i ���!R/�b*݇��t��i��2����WUw`y^������F@��o�̎���(G�h��T�5�$�����[60&&f%ikޟV��3��߶� �ϺPߑ��)���:v�6P����X�X;Y���ƭN"�I}��>�<O�����0.~��mw��d^��SG�����	�NO���&��e� �j]��B��l�?[���WQ�Jh�aTXDBOO�w�桏�!c.B�U��mxA�j1*�e7Mח�6	DhL�՟��K�"�V������O����2��ĺ�.F���ז���������h��(=&�y�ԩi)WH(r������9��i�r�5g�yU�0��4��JX��Qm��LSLp��:�$���A?Y��Z��/����� � ���L��Rb]��*��=������(�:�?- �6]�J�N���aY��m2z����]��׈B�i����Ǹ����'�o��~=SS}�~�����u2����SMQ��+�rt��6&,H^�y��&�A��5��f:�s���~&��}|�6YƼ\�_	s������!�^qpՅ�2�ߛ$�g��ч�r}!pQ�����Ǐ�U��>�ᬾ:�C����Q�]�v�Q�V��ZJ,�(� ���$	A($F����Y�s0e#��<��0����n;[[�����C��^���(��^4ѱ���M�Aj�nyc}��\��i�$$\0�y�#�H�����F*��*"Rɮ|�2�O���V!!n;9�C5��ս{ ���
� 
�7���N+��8ȯ����=�TwSI���"��]�	4��idwYȒz���A�"?
�@	G~�h��@��.�)E�h���r�� [��L<�X>�6���3�
R-��=�o�s,�����,~Y"��c��_'�a�l�ޕFe.��4D�o����P6�}�� �{KS����/�(���:s��ܾ�kC����y�'#�ϋ�W�Kr��p�����+�Bx<^��n��{�l�1BSx�6�Hx
���c�W�B`�#p�Y���������۴�ѽ)�!����+��C����߿k*�"pC�3�?�H��!�0�eh@�Qʣ�)��q�@�pHv#c�����o���gW�f�rws�	fH���ꄈ��� ������7����.c{(���S��2�3���������仵�!M��;J��[&ͷʪ�S��"�|W��gk97!�!%��,��S�V�0�����u�8������5�2��S}�mv�W��#~�H�
:���;7E!pf�lQ�>Um��(�^++�v�;���Gl��A/��
c,M 8��To�3������};#ߍ^�P����800�Sh�������1�0� ���-�D�2i�
���S/����(f1�n�2]��S	X�O�5Zr�y	��Eԏ��6]�� 9�w�5�����>n�y��?���wa,g:::d2�X�= �	q�&=T���y��r�:�m&��ŎPe�y�h!Fۋ�*���h�:�����ĕÈ(����3��"Ku�6�9xz.p�R���,�i�����N����J�MT$,X�
���{��(�0w¼(1�C�I/$�|�s=sh���zA�L%�'j�&�Hu��y�%��)�9\_}�I�=3��?�0��_͎�����������>�Uٛ�=����@`^���^Kcy ������r�c�)�h'�]b��E>ݤ�E���BE�K$���C��S;�U��Q�s��m�D҃1L�z�w��ڟ�Nz���Gv.S�������'OP`&N��d��������_��4v�w�����@��h����Q��g $>�M�L(�$\�䞩A[>st?�MaqqV�u��-$%������_�?/�|Na�)W���~w\z�+Bl�GC�[K�I+�����O�#���V����^L/j3�*	NA��w`^�G�~L�S�C���\��k:���Ǐ�m��������B�pi��t���͎A�a!ϼ*9@�BK�	2�i܍��4�*�,�Hqիq���(�)�d��kH{��M�8@�G�D��!��>m.���F�1����x���d��4}��_SUm�%6&���q�(���Pgzp�m����|l/�~�yݕ�nj��Z��۸םP���3��%�|h>���\��aFI)<)mwQ4��%���MM�4H�t���^.�!���I7��E}4��#���G#"�BȒ|殀E4/`��:b>�`���h:����nVXH���C�~�ۍ�,DDF�z���A)C��9��&w`!���M���~�d+T<�[�Ȫ?1|�}�+K7{��$�&������I����/�Ss�&�w�Do��g��@X�*SE���'���RP�`hb�����A@��M�����ׁa�*�L���hw�0h	9ũ��8���ϟ?O���G�K<Su�����(p�����OB,Q9�tKDRc&�"��|�p�����;THi�=��I��8+h����R�����X{)~�Bu�,�;Fi� uj��#Id��h"����I\h&�_�%�(t���튵�xt*�����(�/@����9�?_�I���,��0���K�f��y~���(�>���˶� ~w=G<g��<3r�b,`f��V�雛����������}�����S�!�C�p��TU�@��q�s26�v#��sCCC�!:LN�WQ#:у�	�\D ���`���|dǸ8!b�9w���~���fv����۬��~L�}R�{�=�<�� ܨCbvO��:]�O`�n���^=��.�NSd�Q�AْqW��wM'��8�����-'o> �`�-o��A������z@���X��$��K���`�*]�Ɉ����it�fF�
R��z���:���o����.�ڷĶT%:�ɥ�%�$)5��S�+���=���CJc�U��;1�F�C�NI����N���@q���tk B��^F�	>]���)�51aè�80�E�)�@��0P|���QJ�缓�� 9]	�@5Jooo����ݔz���[͎�!忳Gn|�����9�*g5�k.K��_�8�_��;���t�$/�A�*���e��Ԩ��(0�(ө��AU]#�ٲ��0�7�����s�B�����$��;J����j��.s;�P�慵H�=��S:�KAM�@��6a!��xt^�K oo�3��d�#K�	��O�����-Ӧ�6��)z�]~�JZ�<�S8�J��.+�����Ke�Hz%����R���X�/�)Y�х��C�O��(E{���p��5���
A+�����.�, ����ܮa?-�+�Y���6�_�7�o�����x��ET�>ú%АЬ_U��`|<˼/jUK�I'��vX�ȨP����ǩO�Hp=����v_�ň�L�A9��V�F?G2�ܚَ�ɽ�M�P�l�R.��J�	�ǃZ%��tg @�d�L/z��� Z5�%'�Y�N�_ؒU��E�$e��c|� lG~!�^1,�BVx0m�m�U�!c��d������&_��gw)�p����OqПB�V�Da|��P����@���@A�BI6d����D]w<����R*Z2:G	��7-��+�"#3��4�8eEY��#3���AVV2K�CH٢�u=���������<�}�������r�H��qj~���^����4q�5�]U?�3g�{T �n�H��(���ь�E�f'N&�V	��䳟,�2�s~�OE�H�mv��N�#�]�)�O
Ͻ��u��o�44d���I/:��vA|�Ky-��yT��29B��'�<�?�X$B�W�9��MN�5���3�goU:�Ci�.���'����� *�Tw�g���͟���R����9����AT@�����E>����χ;昗̌���ŧ�p�!���,H�#R���3�57[o�����n��`�	�9��#�u����HC�=���B����V4հ�����W�'˦^{����a�>[���s���'Mu�+p�y<^}3�~�_�<��C����-�o�&��ާOYԁ2ȫ�ޒ�x�������ߟ����7333��}�Ŝ��2rM�)�W���(=KW�w��������`p��}����^Å�ɺ:S7���nF0��,.v�:�竿-���� ��F�}6K7�M�>�s2���U��:j@K�R��+�8{�UU��3��?. 9���s�b�?�0����#t�	���1^|ݧ�����=�'�6��ĩ4777�6t ��"U�ysfrO3�+�N��x��<����1W#��;��R��������Z�a���|˞��� �#$ԩyF�������;A�蝚�ITz|�D�\}�[�KKŗ��aZ�Lr� K�'���4��;��%���qL+����~��+X�����6%�����x�knf<���P��
zl)�M)����!|��b�ۘl��w��ƃ�v��3O/�;d�4�`��Ţ�MI��}B S� �	��]�_qk�a�����ի,K�H��dEQ����B��ƽd��wߣ;.�B x��$G�̛�
;��bp��M6��UE�HD�e󿗓���K���T�L�ϭA�P�\��+ɱXs�A��B����O��ZUc�<	|Ƶ�w;�Si�r��;ә�D����'��H��+!�@�P9�#z��
3IlP�&\O �`{��`������O�p�ql�*���&��Ig��ܣ��ǚ]6[�;R6hK��@Lk�Ҿ�����K�߬��<O)��8~�v��H��Oj�F���{'����b����ur��}�P��C����u"w�c}B��XK]]��u��p�κ3����NZ��qiiV����}�rɽ*4DP�> �GT�U���Dh��; ��l��U�T�������8���ώ�����\i��d�BdI��-߃���0{;���)sP�ٯa�O�VB{h���GX����K������O�+Wv�!OxE�{�����d���c|~�u�M���/��q@M8�x���ߟ�Nc�e۲e��e`PyO�ec���}�H���K�	��

�}6�?	�_$ ��2�L�<��!���ܘ�]�����0��4��t��s�͋c�����z�M�.�s�9�R����q�=8�!��A�m�j�e��(iZ)���S)�k�!���f%w�-�f���S�{FGF��#�5y������X��FV�`rτ<��s�m�$n�<]�{i�,�������O�B��mp�|S�w@w@(q�S����*v��^�e����qg���g���p�,Dl}���J�Ӏg\�����y�6��f·��gB��ix���'���/'�G=Ex��a$�	h[��;�L���}�m)7sxx8��k+�-Ɓ�&�d�������zs��'�B+gI�9E�8ᖙ��:&��@�0C���.N�痯���6A,"[J���9��S'��k9��jt+�gO�T����x���b���j6A8�"�|-�+]L;̉���}��!�4���}��0w5ٕ��������Mϻ��,|��gk��Iy%Ƞ���G�[��b�.gg
�YK�Vb4�%�\�p�H��c��#�[� 2XP]$�YK��m&,ȥ��(����sf��Bޔ�m�����{H�Vn?ZKz�'%Q�^�Or�s�\נ�^�hhh�J��[qX�����'��Ӗ���~�}�p"3�Zjg5�p�c�����4�:��1���tN�_rp8�Zp��Z|s�����~X�D�b��vO�E��NLNZ:��h0�2M�ڵ\��X�Z:��qq��������Q�/|�����O0���Λ�Lȝ��e��)�~ZZڱ�e ��aN�Y���(\*{��@��,�,[��O��n��*��ej�?_��Z��[�0�++�
��
�����i�y��s���Vс)��˗��¿��'"���e���67��`�X���'Q�t�S-�}�O~s���������)��堡�s~�ù��utV�+]h��jPt����Єi����ە�=OC9�.tQγ;�H��G��sN�r�S����#��ݻ�k!"�jwQ�����3 t$���N�r�[Vr�G�.y�o��o�������Y��;���Z�W~�J�똾	b�Lf�����22����ѝ�;�*Ŏ��[����ݫBI�-�1(xk���K$_�!���X/�gɺq<��� �],�*1G�?}��F`{�xˌ/y�w+��5ڮ>��7�8	<<ww?���Z��N���3mj�b�*�[:���/m�wL{xQG���!���6�}�[� �����P�-|����!��{�/��|��3>}}}vǷ����Go��������.�5u+�\<a�bƶ�v��o�33���B�y�W�ד`������ߺEs�ܸ3h�Fbݻ";��V&S�鳍��Y��s��x뜕��c�9����(��[ �u�
�l��c�ѝ�4Ǿ}�Ԃ<Ddj��k���&Z~r����A�zIY�kv�Klz��N���	�w@R����}+�k;q@��w��l��;^ʫW��!����$��k�m�*: �[]d�7���x��p>�<�	C�S	`�D�si���QRY����#/(CNI��w`��B���a!q��U�f:uI�7�֭[I4�$�W�6{B(Se5���5f̠���z���exт���x �9�g����6��B ��3���V���=�ύ&�<�.N�]�D���-Wq��[�f8�ZI�����l��k��Ʈ�lI���ר`�+!���};΄5o�\G�=�ϩ���gg��,���~X2����=whrI��qP,�\g��LԨ�-k�U�� ��ir�_�9� � LQ�%N��FJ��o��t��N?���	�s��`����Fr��3G1��)���Z@���qbʠ�T����"a!!�3���U��ܟ*K��n	 Xw�����������,�����M��ŎS��" "3,�Y��7ú���N���ѝJ��>�T�wbQ��������`<~@�j;q�l#����K��>lI���6���qq��eɗڿ�\�}�ca��N���++#�P�ڣ��YNݧ��{�/�s���'����mֵO�Δ�)G���C�Zu��`�z�,����fd�S�8Q(Nٗl�x��$;K=����jo��S�#��'�#�9$3 ��Z֥/.֥w�8�^�)�sU��W���u_�`��63�F-�G-����'--�����·]��r�%�はT�0���z.z����~�4Y��]�
��#����bv�9���]���[�v�n�4��v�j��W��cL��<�6�px �]��}d�xU_>�ć����	�=�����dn&����[�K0�|�U�C�v�K#�!���*�iڊ�� a׆hvR���թ�6e2�i��Ū�����[�#\YY!G�G�!۸\Y����uv����5.@Z�ͨ��@��@��@�k�-!�W�$����˓��ʁd���:��M���H���L{~*�LB�qg�������2��C�;���w�{�u'l�Q�,,��e�C�+AII[�SƇB�~���`�vG �"�	i���<	�����G�_K��b~�34=nA�{�J-���P�ٰ�����|���"s+(t��={
KJ�``����`+K�߃ �4�:��QWGG��d�	Gh���Y|p
����-z����>��dK���p�n=�`�ڂ��Kmq��m��n�Z@�}��� ������^@J9T8�
�OE�{�$�w�#1kdd�X0u��R����tOQ� ��xf!#6��mG�[Wc�r7�:9;�/����������D��rsh����e�x�X����=�`��8v_T����p�UT5� ��P_�8$���>� ,}TUƊ�n,�=>�g2T��!��/zU��eV�r7� �u�FӮ��)FrۡuD�A��������%��9����ީ�[gkr56
����XX	f��@֜�ȽL	fM�ґfP�{a�?�}��e�#x68q��� )�չ�-A����P������W�^I$C����m���������j;CB
�x�+**�#�Cb��K,=A8�A��cx;Y�S^V����؟o��,�l�XC��t�Km�*��r[���_��WN�')�/��~��hCɹ�ga�bfMLKNI�]]����c���Q,��~��0�O�m'�o��8|;gi������*9��y��"5�{{�۸��{zr�Ӏ�I{�=nq��1�»zfg���_�謬�{<e[whg ]��h�6Q���p��c�)CɗP���@���]���:Y{�҃����K' �'0��8�e��Bݤ2��!���V����p�����q���0�N._���4����p%�ޮ[�t�"����f3LW���k>���5-�����౸x D�j
��,�6��bW�m!���R>Pq�E2�_�s�̋w�g� �2��R<�s~��@Zee%�u�ǆ0�[E�}6�Av�]�J[Z��s��X����e��w�0G�H�T�K�^�����1�iPJ}����_d�NN�ǵqS�֥ٶ�*W{|K�",�M���l4��Ş"���bUVWw�{�?�ȾO���u�Ư��BtW�vt���4��H���{�F	a�%x�k��@������1�E�E@��'w^�a!=��#�.rbQ��ǈW�bkw�����]��KK�	pO`�ڇ�����'q���ko���X�����xy<��9�Y�ƥF�x	EzN�|�GpE�]��l�K��aPMgg�\����c�<�>�Ɠx�,J����Yf9sl|~j�����`��G��(�Dis1�����
��drg�\�'�K��-���<uLZ[w�S%��D�4ߝ�훈R��T��LK|�A�ȗ���`	avT�w�0��6SJ�XyOͧ﴿� ���	��]��?����Dp��W��8݋�c�v�X�l��o80/�9��~P42�n�"�#�#�ٵXh���I��NNNe���D��k�<��a�Z�འΨ����w���U���s��C�b�����ȑ�g�+��l:֙uA���`O9��;������I�]�T����뫿�K3فq�W��Eü���_`�P!�Sz�J(��_��瞈����Q}��w�}�K��Y`��S9׀���s�!�:��kѠ������l����+}��+ l�*#d����go���^̸m����0P���L�~h����xw��1{`m����D
�7; `3��$��r�>�����}[��Y	���'� ��T����b�������
���!eq6t����%�B�Eo���!G>o�&p�����2`��j)m,��)��{ڨ3
�,R���}P���2qz����5(�.ӛ��㺮+�j��� ?H]��W� �xSd��F���Q��U Y~? 3AK��� �R��2<��=��k䆱��������٭X�
���`�r�����{;�&�4���C�e������<{᳇�襝1'�,��-��W*�\�s@N���l|��ꭠ@W�Fs�k��"u�
����<����Sa`�J�zoD�+��Q@�3�V?�]���
bR7��3����5P�iv���l�Q�Ux�+�!˴��e��������N��p@���,���oxu������\�U!�m�ȣ���.Qخ{f���c?��K9��I�e�:^��+I�����?N,����b3x~!"i�"
��mS8�2dX`����XpbO��8V �����R��eъ߫� C^ee� ��?��,����h���%���w�]mm��;�2l�F���$�h��ao�ʛKԔ�����W�dWBWǫV�D���ΪIM����9�g0Vޞ�����,9�I�eO���:�w�#�$��\�����u���M#ȑe� ]|Ss��XGFٍ������k����?й%�YO����*AR`�-�~�� ����.������.`�}Yq���_��A��6��d�Vecc�߿�gbS�/�j�7~=�P{��0hz�	��������e"���U��4��� T׶��Ȏ*����ϔ�|�kH�<�M�di!�T�'�<�X]Y�y� ���o�h�>ot�F(8�e��(I�ܘf�ꨓ�ک؛��b �����GB��I��7��^�����OK��pŤ�)cJd)NB'N�h���9+�VLK�!�S��+�9C[��è\���~FC�B�ڦ��X
@2 zO�"���)�`V��7��C#�WQ8^?��W�8?�B���EYʜ`�}�ů�tObbN-p@�'F�I�y�x�3;c��.�^�;�xk�6>Q��R�c���w�����޼�C��]�H&ss��g5��-�ݚc����n"�����#��B@�+m��L z`ި3�D����%��ɀDŶS��`��A�,�1"�?ŷ�Hd�;��I��`����5�8�{���Z�΀��}�y�>W�1�����	-���@�g܁t�lQ�g``}�%� �F���hY��kk�'��{��[�� ��j2~��[&�<Z���L!�����o'�9<nE0O~mML��7:[�
�c���s'%5��k:74?�C!>�Ҫ�����&u����ɾ}�V�w��
�u+��C;?Vx���1�Z=�uD�q��P��㘘�5/
���������㍄o���2�t.9�'�a���#�ED,��6h�<1��Js����"�m@%�Uc��%n;y���A�6� Z����^~���x���)9@�|iy����\�SP�)�w��$�
�~s����Ά�m�\��P�*�RRW%N)}_j�K����ۇ�?E����B؜S7��6
���,���v_�����f���}�(�h{��F��P�57/_S��1iNQ���g��"Z�Ņ�b�%�Z#����?>�hd�S?�|��^:66f�flh(fx����R��	Í!���]gY I���]v�=�x�7H���bgҨ�֝��I����G���Y@@݆Uɤ��{|�/+���RS U���Nz��FK=����!��V �y��e	y%�­�@��ݡ×{�f��M�5| ij�nm"vL���v�p]"�19ie�4u.`��N��E�l5��tŃ�bB5^yoa���
������gk����5�v=���Jd��(����!�3��<�h��M����Ap���`�| �y��Oeff�QX����re�A��g��Q��'DD�/�Y���w�?��cQ����RX���OI�u1W�X��ٙ��@xT��~N����t8� ��G(� 浐KF�[�`pf��D��J;x���\����9�g�����2-$uV�\�'����.t��39<����.��i���4��w�rJ���5�\��5�`RC�d�����Gwh��]
����j�sv���u0��	WL��GHT48�Z`	SL����0`fc��[�A(g%���N�51)���i��pE��O��=O/�x�W����u��?�@K)|���w�ը+�9�c�e����R+�G���#�]F�VĊ}��(K+EX�����gfg�����t_���X�n��9 =gߊ��g�WF�B�3hl ���F��>�������j0�Uu=!G�uÏQ�W� ����KsN �*.��y��n�9�:^ٍ��$��F14�	��j`��`�=X(�';���w�់�#EJ�|�3����]BhW����!�mP�k)���-\\��4�\��uο����̟	�ź�w�,���~��V����G�4($��ǧ4{���lbkz�^�����Y�rt	B�+��:��'n�O���f([KK��Ӛ��AZ����^�2��Ń��d��(�����ۿ~M]�9r��@�>}B��B�5�I��y+�\����=W�nw���\�,�ԙ��T�v7� ��[�N�z�C��W�X5�gP����G
7�V�x!b�Q���a�@p�)V:C���d���B����B�v"�� BBB���?Ä��a������B��W�Rd��~��@��c��p���⟁� ���I>a��nۙy�5q�8�ܩ�'O�޼�[��j�[?����@M�[�c1Еٛ��'������ |�P��.�r0�S�Rb�q*p���3�Y$'�� _ߢ?�e۲��<$4��`���� ���I٭,͒KD���!�� ��Lu�1��=�iRa(��-U��;R����FŴ�i���&|;�I���ݣ��M
=�㘟�P=�~��)��";��v����Υ� 8�-̬�:$9�����k>����4<��4BC,�C=�E����OFD:h��!o)aQ�+����1�G9�����p`oӴR�.����`�8:�="N2�����u���-q�M��U�9�
0���	��~}\F�> �l,"����iqhDG��G����.�,�|������R�Ǐ��;�Q-��2�n2ȡ5a+Jl�#���;~qϞ=.@3ԪV9C�[t�ev 	=��i���Bwu$�q��s�.�C����>m���6�׋�λ�>KԵ� 6ZЄLBmK�]ݎ��i��*�} �5�g�b*��:��t��ʧB��3Hs��pC(+ӈ\Ay�6����.�]5�վ �"_��g�a�ll�=�L|΢�W�,p9CPX��?�ELL{��`^���8p����u���P�R��,�2�^�r����AD��Q�$,�A���W�5J�N��tF�mhd$Ěd3��s��Gak�m�"6� ���$�'�a̠�Е�0�'���}4_(v����YB0���@jY]���6����f����ˏL}��S�|���i�]J�e�S��)=vgH�ٸ���+Wc��J�{�a��յ���b�{����L��H0�r�_��cĜ^�lU�l�0�è��񉨴iQ���CU� 4\�w��8���DO����?��Y
�,Fݨ���\3	����O��]SS]@���8	�����`�<�u��?mv�¹y�����m�;F��ߦC=E���Ie7�g��J�]t�� ���MZx~E���W{:��j<y	93�%뎆�}���K:Lj�,����kJ�q<<��x.K�����^}]�꣤�D��R)�7{]�6#0Yo ;;�%m\������V_4nJw��L2h�rAx�{@�c=>o&+>!f�=��������fȻ�V�;�y�f�l!|���R���jHĈ���P4pϞ��M��X�4tK%�Q)6=�8��* =5D��6�P����wuWA�L����2~�������/���r�5�n ���g!���l#|��`��ʁ���l��쓸�.�I�M�a��{Y7-8���M����Jf�V���M��h����@�W��t�Ѽ��q����^^�:�!/�|��$]���MM%��0Ei3A�$��CĤv��*�QTTt/k��;��,F�8PG���L����X-�HicU�8.#���wb-+�X|���]���}%���hc?�y�����k���4�P��g��m � HH�n,�U�̬(��t^k����L
O���ȃ���GS �/���&}�؞�]�<5��<��y ��q�Z�4��+u�B&�X��� ����y^Ծ�\L�i�����5ۼcBl������w�
�t@�jK���2���5�gkn~o�@��Q:�s�۷0;ѹ��]��d��]�`��P�?	�ք�$I^��.>"�E�^�r���*���Q���I�Q̊�j!x������P����gD�tg~��9�*��P5q�X&�(p>�ʟk=3�2�y���b��xd��\:vbbbT��dp���ACT�yt�'�6 E�6*}����@��$��8hV?����mЦ�������#I��3l��k1��GMܖ�o�� ��V�|������GP9 jo�T!,���	������ADT�R#�$���_�2m��3�,\c�N��{����}�'\�A[��S	Wŕ����@��E ���2.���7�v���:�G�*J�36#?�s}��;�,.�,=������di���!�$��>]��qÙE�ؾ���/�Av[�N�R���~�fߝvy~���ObPak0yF���ާ����2�o��%���.�p���ڳ(B2鶶���wf�a��9/��$)vuk�nln��"�Z���a����8*�Hy�T�bJ e��ks33__�mQ���u�! ��:�ׅ6<m'��]���E&|G���.]�T�\t�T��ASAA��a.8���ҫ4�y3��&�� ���B�W��9�����x�]��nSQS{��7���;�e8C[�{���*�g�I�<��)s��ߝI��!_�,e�+'c-�^H����4�,D�;�2\���2~����LͲ#���4���28�E-�F���<& �?o���5����е��	p_���O���8���M�)R';47�����䊣��l�$c�t�!����= I�)�$X2���0�;;��W�w�&B�v��)ΝB+�5�r���
�c���r�e }�'+؝fڛ����w�
���R��6�?O�w�̅��ƍѫ��1y�"-g{�5k�u�YK�!��z0�j�vp�����W�bwO��Eb�N�E�>�@f11�Z=�0�U\���:9���%�Y����d4��|c�����> 02�pbg��H�� Z��<t��!!�nw��,NT�T�O`p���/��J{GG���FGcw��N�A�r:�|L��KMIQ�����ؐ�2�n?�9:���8�G�W��
�1��M���w6����{�MO�������,�+MV�Lނ�o����e`  W��
���	`���{�v�EGE�� �������@�g�ms�ﴲ��I?��i�BO/Y0�!]�y��z߃�,
�*��W�4l"��%$%���V ��D�N ��A\s����e������������8����5W�Ϟ�>�|.�Z ����Ԥ�ȸ�I��%�/�����5 	�>�x�zvSSSD���ÞM*
4�t&YѰ��ޘ,�@�7���^G�]4F���Er�G�IC=�Q.��� .�K��b&���e�������mC��m<Qdw�I#@�q&;��\ ��
<r���G�ؠ��-�I�g������|�:���XF�2���lr�)16�p����q�^�_1�^��ZF� $���9Z���H@�+�",G㚋۳ݨ�5�9��p��� J�P�|���ڽ�$Fấ�_p���&�0`�,�����B)i�1����}�ʜ�}S>zX��D �Ac*L=w�v}H���^��/^�������8���<`Ow���
����k�EE"�Ѕ?��}@����sR+�\ª���4N�Иm ��Y�/}��l��"�|�Ul �pG��D�t�J�����;lF{��(���w'<�I�\����ZGccc#��!d�5�8YԨ�܈5�2�`䅸�{bŉ�y�s��|zPHTl�ܷ������iF������Ly�X@:�-�S�ÂMw�D�'+~6I�,�Y@��.���9s+5A�@����һ�\Tq�ӠiKY�^]���}������=":���4r�uBBl��1,蝋D�ЈU��|^V/}r��g�vT4[!�Z�
�8��-�zđ�b��[Z��; .-R\ws	:tx�f��_M��	1&zk} s��Uڷ���h�B���=�K��]r�#�p�����U����R�ό�Ɣ���Lq�����|l�E��O�`0����F6 Ԍ�K$M�*��p�C�+�"��E�V�.O ]-�W-K�f6�NKJ�Ly8�T�Y�n����J�G���E��d����Z�&$�U������x��ߒ/�=i«����Ǘ��Ez�����������?��q�YU��O�]a�)���%�é�+��/t���-�^	0s���c�c�ck�ݵ\߈���v�o��\�Q�s�������JH���(������o���9�K鸻 vkT,�֢�g��W���ko�p�t*�o�V���f�J�=��3��ZZZ�FO#��w��T@�s�O��0��w@�i����vw/�T2Z?�%p�1�" EZ�g�2q]Ǫ2�i8ҁ�q.$Y���R5�#�ľU(��73����}�7�S�Q�H�/���<?V��څ�7�95��@ɔPw�;u-(�5�ܡ��Α�Gϊ��ȜS���� �i���L�[Ǳ��۠�Q��Do'�W�f���uqqRa����۬��NDXX/�M,uWZ`0�Z7Ui�;��0 3А"��G����6��)5J��S� *Sc�?��Z8:R0� � �Qt!���[62c�[z����aN,��z�����Fqع��izwQ�v��7�?�$)E�5��jWA��U?��Ɨ��s��(�����l�Tv������`
���B��B����r̡��C__�R$?7��k��"�^SL��TEJ�OO�Y��b���r�
A�0���ƨ`M\X��r�Os	ž�9�������7�\���8����Di�GB� �=3S8��2�2dck��orJ��V��u[�Jr"��;�u7����K�4y��l��z]Xxkbj=���Ւ4�Ӭ�Y( �E�����I�����\`4��=�y�0��T�b����;���eθ^�;�q�Kr�x���	�Q,cj?�3�+\�;Jyin*eu������<ٷ��Z��͛U&��X�唻.<&�}�c޶tÂ����w��'ԙ\6��<]ҽ���*��BXğ�+-<ZN����E�{S٬Pn��ONI��y�x�"���c#�8�"ޫ�G2Jy�sm �V�n
���}�즎����xE��W:%[��~~o�v,d���~�7Ԕ8]�wkxP��i,V��)�����Օ���h,��v��)^t��q��Dq�`-��g׃�a�u_"���H�>zE���� �A�r���� t?�MO��g_OQ8��pF�b�J�� x��rC,7%<������j����v�1~���ڗ�#����ϵn �²�S�*A�M�=Zr����@~��stq�$�=(�ܫ��������n�d������,E��O�an�!G���ߗOT<�S�3�_�鄿!���]("#�V����k*�+��
�K�&�K006��&U��NL������l��}$��p�A�f���Gqa2$P_
�4x�E$���SҘ�6��J�d�exg1*�ݵ΄���ۣJs����� �;>��+-ᵐK�v��X YF�m�6rPX3E9y�o�A��J��)�H��n9�^<+vG 6?�\u�	�}5��x�1��h���~4`ϩ�q���}�4N�����������)&�$� W�{h�c�R��?�.J�V�#$�kf{m�i!1�T����aV:������1��M�KJJ�B���_�L��4H������U{Q�s.�����mF%���^Z���Y1�����+�Ҧ�	�������Uвe=7�577O���Tg�ⓣG�YH����%���$ d{\��z�R�5��nFN�X�uJj��*���nŤ���L���d9�z���U��kyՄ�;B�dҶ!\�z�:��[�����a}4iZ�d�ן�{j��{�^�|�����{�;!�̩��޸�4X>h��Ƣ"��\͇������ ۏ�|���a�E���!�B�!b�^Ԩ��f6_C�^��ؚ
��Y+�om�c_�B��-i�k/�c�7�GM[\��/�>g�D;''x���>.�[5��Uzx����H{f'n^@�n;, ⹁���$�O��ٜh�Q��i*.����+���S��u����o�,D>�گr#�zMM���v=6S"��1�������l��l*��Z��o:����/����S������zy� B4�p�O��.���8�]���{7����8c����U�̄��:344�<T=4�7x����!1���7�G}�;�r��n��Q*�<jj�R�3��h@����5Q��J�������x�/-��>����}����=�a?:�;$i�v���ljd�]jT9�h$�˫D�E[Ⱦ(�D�G�;��V��	,������XՈ�O:��y}Έɶ2v_���=��s�k��E�(�Q�$�c�J�󉞁��7�^�������7xA�k:�[c#鮊��hDX��p�#c��������.a���]��bM��<I7���#�}~�?&	���'����W5N&�/	r���f ��Y2x-O�W����ۣ]uQ��z�ͪ�����%���&����J(��W�W�����h���|�-
�ϙ4Q����9EW��a����N|੅g��uE�{�OjW�Sꛧx'+��,F|��Ngh>X�V�r�:9ى=B�.+�LK�a�h�����#�qyb)��";p�����,F�uܪ��W��Qǧ����t��4U���P/�9�S�F=�4�ݥ�&�����xRʌX�M���d�TLy�U-�Ma=�5���֛�-�����kYŝ�ޔ��R�D���E�@X0��=�p��AD�TU�^iz���C�3̺I3NEncd��꯸s�����I��A���H(�.���CSA�{�y�.�b���)�mo���?;�z�Ѧ}�qՑP�P�6��k޽��.�q��Y���-Z��m0=)��&^g�^�0����W����v�ܹ#�:��5�*�pŕtr/�U�qۜ�d5�Żwth�k�#�:2�l����=�(�eX:AT�z �:�+�����E�Iۃ�\�4�\����Ӵ�G�8Ph=��Y��"��^�|Fv��~Y�7�	<F3C7K ��@
o��Օ�c��W��ж�2��CĦ���(�֎�-�D�qM����֖xT/�k�ʖ'�id��z���˷'�>�Z�99�[�Ǐ�ߺE����o�˅�� �X%����Qoʄ�9��Y��CEm�;�����!�2lR�Ak/.����X��}K5_�V �F��J9�ä-����m�nPbF�	���u_�Ķ,͎�Ɗ�1�ub�#��^��y jxc����5e�-L
��:�/]*�Ԯ]��j��$ �:�5�����3_5��<�Ųe5��ǓƱ�~X��=�g>���gI7�,��.��l&��I���x��2|9#�tJ/Ǆ<E�ŤLY�[ɂ���=0Y\L���3���<�DG��,fU|`)U�P(	1��Q�]��mqN<�qcs��#�B0 �;� �+>:��]2��G���7��1ƒ�ʥ��#/i�o%+�j��)yϘ��I���dg�՝�������k�o߾2������E�?R��M�E�'��)��s�"���Ӄ��		D)�Y��G8�>I):.��ǡ*�g&_����)`��y:�M�������e=���y��}-';Ӳ{̞����R�}�E'n���J�8}�������&--�3�Y�w7�:�:�r��և7��ڂ��ڸ�B�asW���&Ԣڋ��%_{�����(lo�N9� 1z�*)�4����Ƶk���.K3�[��� _WSk�\�x�����'���[ø����r����88j�������uxx8?���{1�� 5qJ�NW}��n����[�m��h}��o�c--C`�g��/�\{��O�}�L\���?
c��W�c��:.d|�h(,$d�.�ټ�ޯ��7(�گ�y�(6o��G��tϲ�i�J�'Z�	�I��I=������}w�T���Tn����K��H4�Ѭ���o�c�����y�eUU�o�4ef�.L\��Z����?����u�!B����p��<��Ғ�j�-ԁ+���k��rR�?A�K�g���.�A��rF1��=ک��kcfV��K�G��=��2��������{xYy9$)�,�%��I�[�r��.��$��ލ����n�Y���1u��"v���6�ng�����1�Z�Ѐn؇|���2�q{Ö��(k�1�;%��^2�##6��wG�x��!���ٔ�����S��Z�{|"Z�5����iUQII�u���ivL�}�
5[<�@n¸���Ŏ����K���i[[���{��|ʷhp鶈�>r��(A�LOL�={�8d"@�A��&ݲ96�|\��ʙD�������޿��6FB\����(+3|��~C��������_�?�Aպ�h��lubvO2���/�czj�9J�(+e�K&�_��eT�(j3�9���8))��ʪ���\��U�?�8ʩ��CȢ��͉U蘘d'*����k�g�juN���/3{��1N�tqq1�����O��L�"'?������I�^���$�ƍq̓�[��t�ݭ����w�8�c��2�Z)�y�[}~�T	
6�?���"�%b�p�MOOg
Ԑ�y�u6p�uw�E���d����������2���'z�զ*��a�*��/��}��@��`V[	"+8h'xM{O��4�K����jD��F::<����6j��M�a�W�n�a���ip'���'�]L�%ꍍ�7Fc�]�i�Y}�n��a-$��󡜐��,--�,|7���Ш�e���bb}S�+!�����<7��YX@�D�%�	=#'?�f�8K	��>(ƞ���{�n�?����`�|����\5���L��(��L�y����KB�\��ĸ@��=`�~�ycU�E�0� *�^���qm�������iF}��]w��$'�i�<y˾���%H���6������m�K{���GV�T)���
�Ʒ��*<�m �y}p8ל�-C�l�)$�r�uW���׬�I���9s�d���|+�m�"C��^�����&�]�^1�P�O��ʾ<R��{L��4O�|X��W�P�^��l�3ȿ{':��w���>N�����3�GsR��>�0=���H��7� @�D����wuQh,}͹�����!NDC�4M��4�t��?�r�� P7��G�V�r�_��zI`"���� ��*���۩��ǺTD���̸�k�=j�9�ϐ/����u��s��Onii�d��ϵ����b ��"��W�?��y�����C}�5��\����b���_i;�_\if�S����	������O�xEg����D���CR��y^�xx| </��o~~���z<ȃ��H�#J?�[B���:�H��KAv��T�@�c1���xG�C:��_��Y��,ă2 ��v� �^�5`�X̰jj�Ǻ��+�?�f"��/��`F��f�CD��c�L2$'K�ة�𺏟4��tO���ÉKF�F"�+�����Upf���ک Ӊ��w>t2
/>svvr������� X S_�A��A�SѲ��x�<���N��m�(��+WQ/��U�xM�%oǹ-�OSSg��@���Q\�}^\�ӓ��U"!)���_Ea�g�T*5Z���^��[)KNZ�y�@�|����+.fQ���@�l �%'V���M�߷�o:y�^�Mì:Z��ey��(7w8�ر��,���viD�ۻ;��A�|��&~걩��S�������k)n��u�_��fsn�xC�UQ8���g����E��/<�TU�}��aO����ϕ�����4��avݷ7�Xn\��y����K��wh�iJT!�c]C����.LoNB�9-�eZepƅ������\�̟;&>䝾��3�;���L�I�>�.��x�h-��QW�4�o@d��Mx�B���,._� ��nnE@�̢Թ�ˮN�|���J`���j�~�6�����up�"����	�<}m�]k��GRJ
�.�(ᛀ]�YYu�Gpm�-o��͛7��k��Fp�D?�6b��C@V9�¢���#q_�ۇ ��t�[ׇ�/�/FO�B�D���ᭀ��L5-��4�f�I���O���t�O��:�85kk��w��`
]z�����������}��_F1�9u&E�������:x��L'���_-����X;�m�����^^)[y��iH�`6�5�h���8�,ǯ_o�.ͼ�1ؾ���j����k�z���/{]�>���Ĳy����oQ��z�Վ�kǅ��|�6�A�����D����o�EE3

�����ݛ?X5��*8z���!	��3�AUK+����	|䀒�r��{�jp=y�B� ��6��>����ju��j�p�k���+{|�<�/(_`��>Ӡ@f���_nVT�#������)�"Ɣ���M\��C�=K�dNէ��~y�0������E�ң�;uc��
��)��r�u��!ퟜl}�����6��_��Ǐ3x���<�Wc#�m�����ƍ�A�E)y4���]��an�(@���y?~��V�C�1w�4>y�9o�"���2J�c��8N�?�5� ��H4;n%Ao��}�#���-E!2ʨ(�,�WyJv%#��H�-3[B���"*!���)�EVv��%����o���~����ӣ��}�u�s���뜛��^|
D�\�
'��� 2��oا���K��/�*�B@�>uJ1%%�0�4.����emJ��"RR��/(���a�E	iΟ�C�!�sƀ3w�
Z CUN%�`�gQ����T�}%�x��J�y�S��@`����	D� �����))�uK�ׄ���]QWQfe�I%B��j�v}���%%M���f�s �^|�or��1�T����f��K�5�<���� A�K�bnyO	�� ��^]<߄�Ŀ.�i��T;��[7ݤqV�{��+n2+ne9��;w�y�6�[����~D����jCTm��������N+�v����iO(%N�*�m=m�u�D.9��qG������A�	Pߨ�� /�"�<33s�~yF!v���O8�IGЀ�FP(�,��%p$Ty4)�e|����vO�*��d�zW8u<�Um��}�A"Z�
��q������d��	�[�3/�� �l���5���L?W����#����j��K���GDL��a�-Ve6L4(v
��S��?�?�27�p6�K�yV=�R3*���U�Ό�L`?�:�/�s}���8��ښ^�]����T�,�'�I` ���3|�լ���P�2G��+���������S���P 0��O���hy�tm��x���92}�"?�~��|���;K>�H��.c�<�"$��;2)�����$b�)c9��Ybu�J/3�Id�AVؘ�.����(���<�����$-��W��Y�~f�Ka�e�vf�j>\CwK���:.�(��Z��0C��X�$�WL�-#gg�P�U��!&H�.�k������q�kk��m'���D��pK��M������	
Ȼ8D����.|�
�4��-�d��$��I������0E�}��Y��VgO_���-0f����˞f�a��r��2�uNk�綠L�EȎ�poo2�Չ�)tGͮLVК�>�鎴$c�(`B�Z�x�ZF��ן�����M�55�SuT*�f���
<@��e���n44�\�3����bW
��H>=�j_Pu4�{�g쉫���Z�PQ6��Ы��d2V�I��uĦ��۷����z^�)eL�oͼ��G���=f����!�7i���Q-�D�Y�zGg�V�-�Knp��	��#K(��+�޽{gYə!,�ZA\�ʐ�W��ݻ��eV8��r!/�����6�q�7P�\m��3<�+�(F�$!��*$�Ye=��b����*E`��]9f�@�-%(�}%�2JJ�)iYY����de}G�Dp�h��1��Gg�p<NC]=����������r��q�vA�x�
�
���`e/B�tR2��\�~?��~�)�����}�4G�_�Ġ��/�!9�s]�F�'�[���"�8}Ew���G?Aj�z?x���^f�^\_��l�9�kp�C�y����g2��*ѪK�]B)�<NO5	`�,I��ז�"h���z�ǒTN�蠣�P_Z�B�2mTI�����>t��#����ihi�m��E�-T��:���z(��q���-�w����-{�T766����`Գ��=$]Gܳ�мv���:��ٟw$(���������)���jd{��!���Vm%��ce�r�W
�4��R��,
Cyy�U@?F۟���)�#��Sm;���!�f1�$�Ag
CeT���EJ���s�t���z�u��7�����6/�(y�7�Q�$��\XZvN֥���ƓQ���^06N���G}[mmn��^��>UV�/���z������	_-�:#��q�!�*����~�%:��o�{��%��ի�%(w�5
8���X"�_9��a%����`�v�����×����Yq���ǎ�~+�~.{��ߢ��@2r;oGJ�~fM�hoO; *t�!������ *�X�� �!��_�>}  :�LL	 o1�̂�7�B����8����	�|�|�~A�����p?�ՓPrGDDlG
-�e�Q�%$$�G��'��`Т�"�e�Qt@������1&'v���ٺ�e��m?N�����Ъ3S�{�a�s""S��CijR#5�����]�9�k�x�R,�~	�<��f���[;��67���i�/�v2��uP��� ���!3Ō�o�޽)��}�Y�c�R���Y	ZV��}!����`A��՛�RG�A���1`�O�<QQ����R���6#�7(ܕdwATTNu���a����w�m,���ͭ��2�>sʣ����4�:,:,B1x���[0I�2�3�j੡5%[۬��^<���� �WL�fdh���/&��-�KH�����?=ڪA:�͂w#��᭦���^�s�DO-�arzZ�b[9�;�3)|%{��*l'��\i��.e�O�C޳����f�E�(ׯ_���>xP8�n���
NZi����/=������gRf�`�i�	m��6��ņ@�3�.��^�#��KW)vt�~�x�� �P�!jɸ&�E��@R�g���D�
�J�+���(�}f&
rB�����Ϟ�����&��M������.��EF2�i� 	v���Jb���^�Y*'1�� ���0(��!���~T�v�ǿ�W�%���hY���Y4oݲA��������%�/a���P�*A�=�bFOĂ'���?ރ�i��p�IV(�0~�0t���K�d�J0�yI���I{���mse
�ncc#|��!罄x97T�]^> 0���w��P��o0�g���u��;�s>@'��ѡ�'��f���?C�
Ș��ߡ{&�]�^�A�4���������6�pl3r��B$|��n>r�^�9#��v�����Ǣ��;+���H� u?���?ǧ��Hy�1����E"����,��d����6� r�`7����!a�= ���7���� PĲ2�+�F�O�����l`��{}�(w�擛�j�A�:�ݽnl���6��-�g�����H����	��c�@<���UT���
S7!}�?�����P"5�R&k����|>�58)>4�u����#-d�d�PP@��Pܴs�������F��3;���������n�l}G�4Y�p,�U�Cx0��L�@7#S;��jx���m~��0�X���4�_��oV�	���>�Q��Y�('�LW@#�}K'�<�?��XX�x�9���˂��g2Y.��D8�Ľ��̋���X��3{��xJTT[\\����Y�x�J���%�����5�����|v_\��f���������sݲ����=E�;G4L�w�ݏD.d]ۧ�Y��%�&����)���n��*����Y��L�6� ��Q�bC7�2fF�%&%��x���#� e�����q�>��c��Tztl��(���:��ٳ���	;���+DɆ�{si�eu����{��Ig��d�8q��|����m�^��2�!������	A֪�G�vUp7��xqKQQ12�@G�}C�����	�� ��;Qv�O������{SBf_ݸ�.�e@ME}7�9��,����uuu�LM��L�b\p*�/����O 8���`��(
;���N��д�����R��d�K��b��J�ݾ~Βq�|䯛Læ�ڇ񱱟˞��B�%�2KZj�5��@�
�
_�R{�߂)�/.�8q�kk����9�eKT B�j�͈y��H����n�^��
�2�t��;b�2ٖ��ڮ�S�B	���d�������V_ܘ.,,�d�f�[p�ܹs��V�d���e�q"�y|�.���Ԟ�1m`���x���"Z��% \vYLS�^�k[[[s�ٜ"	..t/�L����\T6��p>�p��+x^Vk[������"�����.�66.�h���s%��}l3��W?�b�\Q�`of\��.ӭ##&m��z^������65�4�Z�*�T�_A��n��JJO�J������������r���Lr���"	q��_|�矪�2���}�1"6�sl����+Ft��ё����d��IN�ԥa{��?+n��.�c�1��²���XNµ�X�µ�|ʶ[��;��nʫ��|ǎ�GM�:b=m�Q�\]��D��יby!��On,�u߾�����;.����N��wk�D��*�:vl�W}밐��~N���}-����n��L78��"̺��` 2���؏�>	N��dc�q�s�	�:GF#G,m��A�0����bb>ظ�klԼt�oݣ��qa�ۋ��������Sء�=�ժ��b/���VWyK���R�W�ؗ1��Q����>H�7I�n���'0{C
L{�h:��#T�heK]�"�����'�b�N.������~�4�%�`�q��W4Y�t��ޑλ����?�>9�ƞ&(��mpW����4xKe|׾�v,v��N@��h�D�W�+P���/��_R������P.�l�r����t��Ü?��P�D�i=��v�9�!(�1(32>ކ$�4SM#D���wx{�T�6�(�>�����km�RSшD!'�>|��M�q���h�N}:�Ԓk�&���G��p��#�\��޿���IA����J�����2+������gsF��Z�vq)J4��u�N��\����dʼ,%3�����6����7�},��sz������G�>�9f�c󡓹�� �����ˆ�b�Wc/"o���5B�����B��E'0 [g�$����P�^`��2
?�j��w�A�+n�[ �#z�M~��!ֆs�x��� f!���q�O�P��b��{3�d�a��{��#��5�x�%��x���4����C�y�%%$�����(M 3<�{��a�̫W��-�����o}!�C�~LRY�Ayb�o��*p�?~��7���'�-^niy:55�[\#X\�a�gEBA�`K�O�t:���-���xf�����+j���呋J��a���f0褞s��J��Dv���[lQ��͍S@������{�R�TcL�����v/�<�|~���Xӫ��Yd��<��5Fg4��t�EO��a4�i�ṗ��W��;
2]Tb��at��Q��=���0:t�H[y����(��9^�ɥ�ͯ�t��o;P�xqDgb���Ǐwqql`����YY��y)x{�Z>`�ޡ��j��ü���{3뛛�!������\�NЍ�[޵�9��GJ�@y{㛓��`Xy�+n��R���2蕹m�!>z���v�8n��e�d0�ρ�>���� 4?��gŹa�������e{���1N�'{:??�ЁZD�p#0Y�����WR��~k�3��ɓ����"�q��}�xMWu��zd2Z��>�RGDGߕ��_%�ֲ��P\#� w�{J��
��yE�(�\{���!*;�s��-�ev=9�(��0HQ3u?��� xhd�}C^6��leU�W�_��8g��R����ˢ��}9�v�?���@EE�
�k���2��
������:�it>ff^? ��<�%�rJڻ&&_Z����Ol�2��{�@���/_���1����JvaA����c�
+1R���$��#�YXF>�������`$�KS�2/��ؔMvߘ������\��9k�+#��;�|S��e�d��!��2�hȬ��a0�Dgz_T�<T���Z�~�������2��f�!M�2v�NN^�q�E�q���U����*XA��	 �R��!�΢_Oxxهg�����X���و��-��U_���[�8�gk�MBb��n2�����U]__ߺ��|������b�
�:)'Gcii	�㟱Ɯ���h�&��Q��@צ6���4�@�5ra�un�~s��N�w	����ԇ�<� �����ۙ��r\;]k���@U��H�,������~��]=�\ S�B�Oϻ?�`���Zs���َpvpxq��*jj��<�ma��)�x���پ�Nx������{SS]����l@��rG_;LwܐQ�O�>��^�t�IX��K�t #B�5� g)���5��`j�����]�q�6$�V�x2J�!��c\C���|}͙��k}BBm���0zF��-�b�#C�_�u_sl��]{;e.*6�r�y7��|)��4��[�Ab��͌.N�ݳ�"�P���������s���F���8d��#�ݻ�� 	*'����GPUɊXbb�i�|7���� Y����_C��X���S}Ħ��Cģ�b��M����ee�v�[�QY�������Co�\P�l��tN�/j���K�z2M� �^K������H���|� ����ofٕy\'2� �%���5O�
;ח��XX�Oʧ�w�̦��H�����S�������Ź*/�bk^� aҋ�$��׃�]�v�Wvr�9Ttl���ֻz�k `�G�e�W�dܧ�����jWWW��'\�	u<&�����Y�`�QµeFe�.�w���[Q�Eo/���n{�&)����#Ҹ`�������������AP���'�W#e���'s�<�*��u�tTP�ϟ?���O���.�p1I{���+nEC~G~�ղ���8��PT֯7��?��f`�W� �`X&�D1[Yv��_}���;�s����N�wT���vB���uܚ��:x����r��َ5ByFXXXAН�+����ubr�t��z�$��(E�^[�^�Et�#D*�*[fለsT�E��y��Ut��z}�c����ˏAώ3�u�א� � TZ4�����{�+�e��Pѣ푌7oΣ������V��e��XvL"�P#*��о���y(;���\}G�g~s�zee�v�6�����k,�{��%�%�����5���o ���#Лم�ǧO�
��2�n�(rpp�Q���Ix�ɔ�����.�?|��B[B��ĉ����5��O��I����5r�vE6Ep�@��A�s���gߦj{� ��n<	|����G�,�z�~�<x�^����,�g��Vk��L4��v�F��inn���"r�i�8�m�"�FY:��%LUUU��l��@��gE���s�4���dL��C՞ �
��I�L9���f]��n:����V�
 +F����}���c�u#�7G��[r���w��X�ʯ�4��j�i�W���G{� �K�y�S�\-�z�<:�'��A;c{�K�u��C.Pӂ�b�-�����<ݩή.��0C�GD�V>�E�8����{�lY� 7n[��ZjZ�UUU�s�w�(Z�+E+Vd�B>���)�+RF��N�����9�/�5v�i~q�Hm��p������Qwb_���}���O�`�'2����g��3�����8�/3A^W�;WL�Y��]�9������}&��uP�i��� ��q"�hFu��U{E����}{+x>��u�����D����6q�OuQ��JΟ�1m|�V�b&,,<���n�}���O�{a��nm6���a�y��v��!�j����kh�5O��"���06|��ym`KF��z���><k��ёT��h͖]�!0�Uu�n�V���oV���,[������I�������_�a�H�|u(�i+w����J�����&�CC���E��jn���JHH�a���:W�]>��Ň�t%�v~���Bw ��%���.��)���`H����^D�W��9P�����ݠ'`kDtoDGK��j���������G#yo�cbb..���G��&n����B�z6`?�����!sO7I�_�IMU����!qx�H<�]M�1���:D�y�2�}����cB8:�(��ё��k�#r��������5��jtR�^��&�����R	�@մW���o�3j�<Z=�0ߩS��Фn��l�Py��"x��=���WTOȑ1귒�2D����
Xؕ�����Dw�~���BI�҂j ��������Bh�DYP-5:�|����;w��m�v��k�6�ܭK��ﰧ����������k8�z!ڃ�Ro����744 0\-dh�-���.e m��&��%!��x�����,�P�~��rL�D�uۯ��V�>��O�Ϭb��rrH�:d���,b���))�Ӷ:���g�QM�(���� &{6�&�Йl�?1���<~d4�%���d�9�9DAN��ހ�B����ze%����@��CTD���k�r��ՕO�顎��lo'(_A��/	>"�.%O2~����r����zzw[[�Z��J���;كe^��b�T��q��(��6�:)Z��g���Ow�ĉO.%0����L��Himm%ESA���aZ�D�F��{��$�������cBBh�I�2���)�v쨁�ƒ�ى} �^�z�=y�۪z���R(--�4_� ��ў�ϟ>�O�R>�ko#�#�Z�Zi�@�N�ަ��_V>��h��HMH��g��*�:���-|��������G7چZ�ږr�7T
��g�K]h%~����KN� 4��;՗���l��Ka���}t��衭���(&���&�񃐯�fT���K��zW�Uޟv0�K���?^WT�4D)h�(�[�+�{p��Ya�M7��`�_�c�w�^@D��<�]h���2pIGǗ���.�<W�=�ݼG*��=�{�'�d;?��>6�+��@�B}	8,dڠ�)�����6Kk%0��Zu��膻��r��B�����~;L��f+�AO����F(�*+*.l�� �xӫ��*т籙�؊�.A�߿����`�����;�.���BVRRZ�-���N1(v�*~��kaȎ����ǒ�Ww<~X��c$�A*:Z�m�6�6"S�5T�
����*�xHJ���"r���p�O߽��U��(��.&&t��͛c��ܓ��=�C�e����_��7��7�cd��cҬ�*�N_���}+%%E7�$ 2��/�551��Tk* j��zk;\�ݽ�;�����W*Mm���w�S��L��ʁm�RhSӤ��C�1��ӌ�n�閱Si��gC�ک������=��"�~ϟӧ�^
�'��6�e?yMz�E^IM�
�u�n��/0�v�<�Ĉ�N�i`�Υ����8c�A�I�s4Ij��IP5��2.t���Pi�� ��*~�� Oz�g{��/�K�K��[:�>�$P���)ET���$��9D�����V�=7Ͱ����P�����g�u���q�>��م���7�_J����ְ�atb�e?��8w����oԗ�.,,�(T�z{��`����B��`c	�V�Q)1㚐v���v�ؙs\�_�JKm}}��<�W�3m���$��<y0�P�=���Ջ��~Ūx����m��m��Or�+�����FL��!�L�<N�ʯ��rW��w��[~��'���*ȃ�h"F��T5��bt��Tk��\&]�+)�9��(�ؗw��h��СCض%mXt�{�
�Nt���������Q*��l�=�&�:����?�����=T��̐��h<�����c�*�S�8Z!�ug��{�Z1��&715�B?	���W�꒢�z(V�B�!Ӑ�K�8�y\��yo�F^�<��"��H���K�#�I�T�r+�$D�h׍�IA�~X��b���q���*��s��-�ܓ������Xt�6F�����r�ťH+�f���{??�6[����m`_[Di�>��������Y�[ VI;LM� 7^�'�%�O��
֡å�,D���i!}i�c��#�hJ@A�8��ܷ�[����|���ut��C�����\M=�+(�sr�Z���.�r�(T��w�i�o��J��3�����Z�i0����92�@�r:��{�S�9}�&���cf�`�Rv�4)���Yt�r��)� +���y���{�n"Dr��5Qy	 �p�$�����D��ڵo�u�M�%Q����	���6ҵ>�ܖ�����{�z�>��:��33�i7r.�
n����� 2��I,� �f�u�������C����1A��H�6��a�{���I	GՖg��_g ;S�'�N�~�R��� �z:�Cz+�N�$�Yx2�ԗ��Hp�Dv�k pRM��ԇ�H7h��SS��9u�rp�;�?H
j	�	����
i>�	1Ɵ9��#t�-V��k���O�E�!��IS�BFY�˄��Λ�����IÆ�;w���Ţ�x��*5�d�Bm^]ת��t߁���9��^��֢�:���
����dϕ�Y��L���՝eE�8�(��)�ڧ�� %ZZLڍ7���ɼ���uj��� �¯RS1p����'�6�+�� ��f��B�ӄ<�2&�T��I..�����(b��I�H{���H��TK�˩������<9��p�W�� 5����-�|����~g�΅�K�A:�G�#�M�@���,v���+�t�S���vN�iI����Y-M�tIV��H�$���b5tD����?�wE1��ŧ,�e��W��=��Ą��B{��~��Z�t��*jj�7R`& uW�s��@l@�i����c���[\
z��7�b�:�f�\�f俎DB�ׯs3�������Y�өo��oM���\o�i^^����9��_���#`�J>�=y��X�|aȚ-V ���wU��`�>�tS}Nw�_\E��r���燹C���gh�g�ET��g��:H>��h���O����ne2�s�i���R@.o����<�Vԑ�>yB�#������9a�~)�W�/��)���G�%:Wc������s%��b�ϝ�,ߜ.��}5�~�_9�!cD'�`&���\X�_G$����ʧ��£�>��	�q;|||�!^IBI�C'.��EӤc˃G����&2~��L��Y"lm �$���>`L��ent;w�������yq�i�J���q���۷Ǔb!�ۯ���q!����ъ�f1O�Q�"i4A�Z膛�'N|4�;?�)�>/���r-333��/y�R�)}�1��_\�Q���و� �hGkE��Ι�r���?f��WmL�o~0�`M��&~}�t��zd$�6�@�����[
�5]�,9��"/:d'���@C��w��!F�������S���a!�6{�t���w��o�7�@;��z���]�������ċ�ʝV�W�4�T�zx��6D�y�pZ��E=�DYT$�4��&�]�wl��iii����v�w�����bB��	M�4nT��{!���Z��2���g�bVOlKVGw����N����Y�W�Ԥ��91"**y}�M��Y_54�c�Z�� �Q�J�:{�)==�,-t�<�G?{h�$�_z*��U��,Yl8�zS{{��r0�+�n�SPP��P��7���_�>=��봕��It��5`g%�u���|՞�YUt⹁�V�{�˿��Q5���Q�E����N����9�{��	)z:a�����u�2+⩆�=�+rfŘ�l�8��$/��Z�,=�q�� w�x;�qצ�c�C�}d��p�On���,�}�[1�F�ib���X��ZP����LC��$��Z���+w1��"�O\�	fdB��l��~˥cOc��Z����*�&�yv���O��{V�d�D�}�U�NLQ��#M����빹'Y���iWGȌ�_˗,BXj�]~
��Bd�.�@��B����x~���R�_�3n�����r�s2r�?л�|�K��&q.? ����U�9r
fvvOho`�UǬ�dxx����b����ff&&�iZ<9��Ja��`_�wH�� 0�qw�U��Ҍ~��e�<��#bU����ПȂ�m�m��j�����'%�����r���
aqO&ە8W�ت�h6϶�(#""��0(�EA�j�d1���������&��z�ׄ�I��\����s�Fv�v�=j���ϛ\����5L��
�l�ե��Pp�GE���n�E��q�'��[�"����W�+���F�z��Z�HH���Е<(4Ԭ�o���]h$ �+5�I�sZ���=�B����0ɬ�3ؿO/ߺ��R3��e�lN����!7�0��.�w��Gk�.Xl!��z�w�_�y�~���V�|��q8�/	�2/!�E�U���{d�[��ƚ2�Ǣ���	���5%�p��^;⽮���|�מZ���"��d'��e&�&�f�l{������ˈ��BbH���wF�"��x`��>FZ�-uq }jn�|���e~r��`����^�N���X�}N�ߞq�w/�Ӟ�;��t�;�u�e\�&��F4�^<W�=Aa{DM-�N���\(���6�kˣ�kirW��K/]*�3��g�Anl�tw�$�0�ɹ��E	9x\�Z�"�����΁2>
�w�r����#��gP�2�Y&���6<���#1�7ݗڷ�7�͏<!�(�{ʡ2Rk3;�[zދ�Tn
Y3Ѭ���5�n6������y<�'��ܝ�O�lK͒Q��RfDĝg�^�޻w:��Q|LY���$P�c�
T���e^��X����u�fi�	@l����5��B-W��v��GD,��E�(7��I$sB���>���S��Y���.}�Uc�x�{��h��M�߿Γ��K��A�?+͞�v=�^�2;h��ޯ�{�-�3V%�Ε���ؾb���t���:�
�:�ڬ�IC�zc}�M&��K��1+.($*�������?�诓扦ğ�Cl`�#_����N�0�!b>�(�#����J��
�u+�������� #j��X�����jD܅�`��ӵ5Jto�E�{��Ģn��o7&�g3�g]�~$1����\��'�bv�<����鏷�e�o�M�m�C����H�cS&!���o�P�*���@Ȅ��TQS���z�r)���+6�ꟐZd��ͣ��>���+�a��k���_��
mUh<�����M���,-iY��;����C<�n��c�W���2H)���f508;`s��CU�q���ZI��EtiE�9���PR*�ɮW"ISF��ihS��<��_l�07�xN~�q"�S[����9��˫���Om��&x��7�t.@�ญ52�Y�tӶ��!�pc�G0�U)1.K�k{֗���ٞ�ڰ�X�El1�{�+�xeJ����\q�"}��mKu5�ރ������Ȯ�����%��q,����m\vk&�}a_������p�� �:84t�w{sb�͗0���&
��=e��z�Q�j��6�͒~q��]w�3q�����������0�b�����gƲ�XD���2[����Ԫ'o������7�"Ⰰe t��3t��J�SY8
k�wb���|\o�Zz��l ���&����r{bBzr-���V�,�K
a`��6#�F���*������tŹL�@jӾ���n�֤"I���R5?ܟN��"���&��#�A�p������:O�4If�� f!���1t��7�|4�IJ�?�\���lU��L�>�23��Gaε�e��`��_�c�?>i��&�<.�v���ea#I��7��(e�{��T�x��?�,�u���Loa�Mr�+��$hCRVCS3�t�g��p�I'�IT���G�	Bןy�;��.��M_�T�`��}�/�6�cW�WtD�sI[ȸ:�dG��⾉��Ƣ���|t}T>�6��.c�gƝ�F�+hi�u,2�ɹo�%W\�6��'���B�9�W.ˬԪS�������G����-���F��F@�]�p��0�����W�[���p��D��v��D4v;�o�;X��C�II�.����D�b�8�����Y�N#��>�8�_�W��m,u�Gy�D	�%���k�n�b(�w�Y�M�/f�W/�[C�������Qm�Q� u�� x�р�(���r��P��(YP����k�߉b�%���o��F��^`�U���ɻE���[�l��]������\��1@ �\߷\�����|&���p���xm�
r灚6uu頟g�(/_dy�`J�BJVk���������1y��+��_� ��F��$�����*7�y�rzB�9N��JRE�mx=�k�̇��mtll`���f��ե+�Q��o]�z�ϢN>�����a��'�AAf��N�Q�ǧ�������DC�w S"8xFG}��'���4�<o�9>ޗ�q,���� ����/��L'�� �g!�=�L��6k���Z���Y�L-��:*���COx6&�7��_��g���ء �>�<���P���,ңW�Nt�:�6K�дt7D���$%u��C���+�q%���_�n^�So�>�_�`�Up3�� �Հ��4I�r�
3��4����DP���N�����jjc���@�
�,�ڵ��]{#���vx���y\6��<�p�h��Rd`�Ǡ��Т���*�$\i�Ԇ��@f���?�u���-�������`w�p���tOWܢ����c���:!ݕ��e�m�B��K�����ܐ���<��=sX�T9|�'�M"�0�D8����i�/����u����[������%m���4^�[�v�	�׽\�^螂㿿�U�������:����4������Gc�_�Y�����䵱�ٮ��[���Y6���W�����~�������������1���׿��;��������E���k��-���i�-�w��M��Fkͻ�l���S{յ)�p�9�$KW���5��?�����7��'��`πϠ������\G�EI�88�e9|_��
��}=���gL�Fk�{��8H��l)����b)s�ɕ����ΊT-e/>\K!����Ѽx�ʍ$Q*��Q�p!)�p_�,PYw�(���,q�3ow�����I��*��}��B�O_|Y�=�+����K�`ei���=_����J������?��Չ4Sr�z�/�	l�^&��\����� jCΒ@VY���gV��Nb?I�^�,��u���e2#��>��^8@z���}����)Z
�����뼥�e�����L/����yK�C�$=�O~Y��MI�P��ȕ}�?ɱb��Ja�7.�>M��$�?t������=k���I�:CK'����%��=s��Od���I���F^�?�s(<�U����]�H:���췿7�ԧ���<ѧ��R$qiD�J��$��t`(0��d�hIZ���6b���$y�h��p�zcH
�2=�C�hP������,w��s>����P��l?��r���!��k�dw�� ɬZ�,��,�KMXS Y�����A��)N��oZ�,;Z@'C`݁蛅�<��%��k�~��e$��/�C��_U8v�������C��_��C��mo���T�ow/ę�������Z���a&�C|�-���<� z�i):C=ׇǉ��-�IV�`P��}��jG����������^�#G�"F���rk��nqK���=�e�O�-jMb1'�{')�O�*1ip@ر����׋�����W��S��3���K�p~�z���Aw�����O�'��i�Gp���&N��m�%�ja�y"ձxV�	G��#��������x�����>B]�LN�Z��1��e�"���IK��8���]T��\p�6�`���f�5x&�tT�ɠ�^nI5�5�-���u�z:����2��H.�K俇}քS����m��r��q����(t�v�����9�����~��Et�LQ&��J�߿���ႲF�bK���o�e����7�_i����:��z_פ��ޞ�Ks2����i\�Ղ�53^wJ��|�q�<��#�?��Kq,�Hh��ᠩ!hj7�)]mq�jU��"�n��	ki/?�6T��=���$�3U��i�W���T��{)��JM���]���G���i;M&�h����ϋ���:*ܪF��s�8H����2y���G���<�@�>z��v��c����d���VI&&O�����D��(��,~�GrR�ߑ��W5�KEq8��p�������4۝�l��ĝ1�����#	��x/<�?���	�k.����k�N�+��p��i
�0�×��#?-2�����J��+J'p��:�泽m����R
�Mjj���b2�lf�@49�<%�z��M�R���ۺ�Ռw�B㗡������Ԍ���B��K��6�}�^�����|fQz�u��ņ�;����p��!m#�=�f��NA+���@8�m_�ѝ ��.J�*Y�8|g�ᅐ� ͖ϖ�4ٙXY7�̔������`�֗T�V��K8f���255�C�jF�S�n�K�.m��MW,.��B6���A�-���E��~O�"�I4���a4N50����Ph��6O7m��N~��E�G���{�n�涾��Lx-��1.�{'�q�c���yh����FVQ�����y��WK��0[j�z�AZd�ͼ��֋557T'Y�RS7��N(�F�ژ��j�;șX`䞫*a��t���e���[.���3�����^��<�n!�͏0��Y))))����;q4�l6�Ax+^b<�nS�6TX�����)������a���t?��N�P;��B�U���u$�Ds���\Fg\%��1}�9���~���e���WܨG���+�4hY����¥��PJ	�u~_���s*\�M�i&R����e7�����b�]���ީ�t�NMu�<��#»!���#I9r}��sz�E��S�zE���~��8A�^��i����~:en+���7&Y�ۧӴ��CBB�x�h| �=�v>�f`�=�#o�O�{hq6Q9*$�m��PǑ�`,ǆ��p{�DD��4���_P����`��=�8��^:V@.�R�0�o���!\_˅��w;ȿQ��*����F\���ef/
]0�@O����|�)DA�0�ѽL������H4v�Mz���4E����j��t!��[9�<	���4��u�A�C#����G���mru�'����TBs��av��#W&�pr[��υ�����t�~Au7�R�������S�b��2�W5r��Q|��k��>����G�f��=�F������Ñ�C�l8�!Z���|z�*�u��L�ꉕA��ٜ��"�%ץunA���E���Oa����j��y�g�)�y畅Q��.�q-�֥e+�л�|������S��z��J�4ۃQ�̦%��q��H�.�/9��T�L��ߏ1p�Z�=q�`����KA�%�����iz����9���Ϛ���k0�6�}�*�}���:���r��a{�f�Xӫ�n�r�-!/^KsI�>�o�L���^�t�up�����G��ev�_����X�����Jt B�2�A��� ��v�A�B����j����e|��6CSS�Z� �vLS�V�N�ӤdeeY��_�P�1�t�	[�,�q�#ӻ��d<%���A~uu�54����_�|;�}�� �^��*��H"�SEȱ�/~/�1m\��,�7�9)�n�n��Y඲`��_�պT�`Ĺ�;U~{����6=�<�G���/�7M���8=p�µ�c]z P����8B�y[�xF��j28�J���dX�bZ�%+;p�zVP�=���U7�^{���Xo�H~jj�1��Il�ҧ3B���CA/����Gz]@x	�K��0�Dj����tO�Z�D�}e'��<�MڥC��d��'zt������m���܍�B#��(n�/\��t���������x�p�_Bk`t����G�8;O̿;hεrUSs��5��aVVi}z�\9�"e/��{��]��k�p��h��/�x.Q۔�*��P�&}�]ȴ�y�ȃ�
��7$d����&��Yt�e��㻛��������S�u@����8_<31���6�iS ;¥����+[��`@H�v���[S�?���ln'�Ę,#
s.ޢ���c`+6�F�U��?��PK   <?X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   <?X@�G��  �  /   images/e086d210-4fa0-4a6d-a74c-91bedc336751.png�5�PNG

   IHDR   d   S   i��A   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  WIDATx��]	x��~gKf&�%� � ���ejdq�"j�kq� ��j��
^T��P�u��^�EY�"��JI !{&��������0YH0�@��|�Lf�m����|_� �0t�h3���=Y_���i���m�M#��4�s������U4nF���!��V =�id9�1-�E��4��V�v3�c�C¼mEy��K"�� B�e���q�F��y<h���&�^�����z:$}d���|�zH! |��� <4g�z%��]"���3<5x^$S���@"��)@��%��S8jw�0ә�:�N�g������A�;�V[3�d��y�K+Rd��C���1�'FF1É�N�e��p:�p�{���AP�=yU:�d2!66��8�t�(>���s耈)2a 8�KJ���q���{޹�((ܑ����jH�����ג��<�n�͂Qc� ��ض��r(Q�L ~�vi��� �_݂���X���I��TTԨ��P]������t�י蛒���geC�y<}ߖ�o��j�f���_��˳?C����`�Y�1OLFj�I�ϢE8���z�^�,4��H 	;H{FF���qǽwchE�wCb[x��R]��N�ҽ��=
C�>�iv:��
ґ#g�톾W/$̛���/+�m�&�j��38Ll_HQ!'+����~���ݿF��_�UR�ڗV&��+��F-qa���}Q S�d	�G��}�(y�(G�g�PQn������`��X���(%fDGG����Ɵ^���� ��u3�޵�L�-����ia�a�Iމ??�>�?'��,�fsOx��A�@�,�y�i���?Ěի�mhM0B�H������w���Сx�S'�7m��ڠ�~�z����cѫ��dF_}��J:��ڒ��6���>�����K �icO�'D,��۶���������W���m�gk�hHd���G��u�t8^���T|�\b'!�k�{�	,�?���F#"��f3v�����t���An��( ���w݅Xb�c��po�M��#P��K�NEjvVā���%&{�{c��p��G�����A@x&��1�>��I�ᣇc�,��	i�={��� ��J�Ŷc�`Է�'�TbP�J*��+�������0E��	6��+���u�\����d��s�o���&?����~؁�(�QT\H���v5��pbF���_�ݷ�p��~ۭ��yFD�N�};�>��Q�5h�9X��1��B2��C�;�h�˫#`����P@��l�	3)�+k1��7�#�	�3%/�r�ˍ	���c���o��˵32���I�{c�;�#�ԟ�,D�mE����ws�u�ĽU>�iRՠ�h�~2���(N��c2 �#�S~��A� �f0��֨6�\�����ܤc������Q}���j��A
�
��:�r��^?(ҷ#��o��ǩttPC-�*��o ����,D�MC���X�J�_�.��OR$���O��j�E�i3圤@�-����qaQ輌��p(:� �|=̥q�F/3u�|����+S0b�>�H��>��ŀ��`0��$�{óyKX{* �x#�,-q�"1�=�U� 2i�@#hͲ���o$PF�v����	yea����<rq������A\��2�������]`�b5�A���k������'N"Ǒɠ#@H��'0�Ĝ�#���%X�ȗ�y��!a�'Ӷ���'���3�q���1�sv���P��t{��	$F������������7���w�|*�gA��W�X�#F�|߽���*h��ڭ�{ֈ�-���i�r`<d�8p�̷w�N��j���XS��R cL����Q4>�7!`0V	)0W��%}i��*T���-����JD� ee���������
��jU��i)� �q���m�/���遇�6����oh|ri�9�F�rs\R����k)�E%RGUU����b1����E�]��눝:��>��c/K�S��b���~BxPz��n�4>��N�"��a~�)��`)��m����9{�@b���jԯ��aW�t�DQ��ó�k�<�0*f�
��r��'-N����s��^+�wZw�f�	< �H!.�}���:��	���X�<�
�q}r
ي]�~�Q��dk�6 v���#��S��MG(�DV��,.<��ޙ'��uW$)"S� �����ͫ��B�e���u�Lx�l��&$ f�x�-Y*`��d23=��)��M�F`�J��p��vy�����O.��U�H�(����קk`_�������L8��v�т�	�_���Yk�^/�1�Eۦ��X���"-�q�g����Z�w{�
9=Zn���M�0q*E����t��Y��TR�>~1D��/L�g�V�n�ѣF�|���_u��pD9�|�$� ��<k�"�=��dۜ�p�Z�G���p=DVD|Q��Q�"��C|~N��\W�,/���F�ZA�%���T��c���-2�] =�%j��Tř�6�/�9����E��[��^Ty:(Hi�P[V.y*����s}�t�2�a��6xSS�����^�C*�1Btj=�-�ȱ'���W�K���6(���/*n\�8T�hu����k74&3��E({�)X_���T��B#sX
q1Ы��=4^�q�ƅ4��$y�+6�#Rp��}�/@�����
$%%A����$��D�O�X�v'��{��ߧ��Q�)=k�!i\O�,p���Ʒʰ�nv�t��M	��0 ���ge�WJɐy�Jv���%�z���E�2�W.�(Z��r导�RTM=d~#H��}��0���]���C((��ك��ރ.6;rJ�;$j����S�&�[��S�ݡ����Ǩ3!t"��N=�&I�
�8����"~�$\���E��i;\`h��zŬٰL����+�^��X@�a��h�l��'K|%j�C�X�hx� S�z����'�����С�f׮Zk�_Ҩ�[�����~� �Y����፞��ER�D���z� �
�s�h���3���e|َ�Qwm؀��݊ď?Fz�y���e����>��Ha8W�Ud~5F��ڸ�I�ds�ə'�1,��!f������`w�b�h�p>+9�,���"�'!��7bI�Gkמ׀�%�V���Wk���9%�S=�a��ٛ#R��/�ƛ�E��u}u��^��C�g�ҝ٧KG�Č8p��͸��[�զM� 7O{>�.W8j��UxL�7��������Ld�w��zH�D(2�y�Å^
���-yb��^L�c�Jt{�=\7jV�[������	T���6W�z�ݱ�W��k�g��CD.��8T :�F=�	�.D�|j=D۰�����o�z�z�=�J��ɖ��G�h6ׄt�k�hh;Q�׵k�����ɬ�I���|J �u�ӳ��yB�W�Y�������3n�,]�.=.?���������C��8 �Ν�u��41�'��
2�����Y����&?�bz��*К/2���g}�]4d�*3ޗ�!:,��1{���F�+QQ�u�5z��bO�3:���77rN䬣bi`M��"�5�rqI=��̎��coT�� ���>����C�SO�|�T҉'(�Νa#�˧τ�{"�X��0@޴}�z�O0�	S��8=`���b�~��D<H f��/�{�K��gB�r/8�nraoH�\Y�=wC߻�h+�3 #!,�7d��jT̙);Z�E,m��	��'
h����G���u��K��W�ܵ�8�|�!�b7�'&��J��A��>^���3QN��>B7�db曭VL��`'ƕ5��@���y�;K	�d�ss ���Я� G��[(��ӢNR���l��t�Ĥ����c�<�n�/p�)�&�Na/��&T���P��䫑0n������Ͻ�Ο}*��E�'�"
�(�.X�jN�E��g{a 0'�{�7��cͰ{���q�����cas#�sf��B��a�^~������]�Q$z�K.�L~��y�-������(7�4�w�/)�s�{�{m1�[��&���|��K3_|�eK��B��e(%P._�.��6o,Z�*0�$��%���LF��Ͼ��'Vs�u��n]�K��;�}��Q��vڟ����rY�*|s`��у�:k� Bk2����8>γi3���2�s^l�2�	��R�I�!*fÖ-Ōy���($�	��ǻ�o�D�<x��p���p���D�I�K?����X��UB�iԾ1K:vL��������U:q�� �W����\��rɛ���" nJ�hT���B]���/��	D��?�Ao�����7IR���(m���N&F=RT���r�b�h��;�nim|���^�@�2�_�~qd�;��"e�=�g��Ū*D/i��KK��$v� ��w��P��)���@�H��<�(I�O�l4�Ȓ��"N�{?��8�	��}�fa�mu�����>q�]i{ϒ
���ݞ�j�R`,1 �8F��;����&�xK�<}9�^�W�~�g��� ������@��3�0h�`���4M7s���0�"��Ñ��(�4g"�t�^$�;�C-�R!O�虩���N<�ܳ�b���b������@h��e��
�D��L��?.E��ݽ��c����x�z�tf�3�B��]Ϟ��j1��"UՐ����!d�G�j�;"��:����E�"~xu5�yyj���lWH5T�^9O��$�[H}}���ȑ#��
g#ƒ���x?�������#�{�m��&H��[zZ�<R}π��B�ˮ���p��O�:x�P_4��G�č9��<\s���kx0B��s�Y<k6��.�z�!� `voނ��-áh�Yl i��h��Mh�!�����$���w�����;.������Ȇ5��>|s�6|s\��cF��8^�a
�M�!�7�'$�oN.����U�q�%��h7������A�؝潸�dP�(,���ųm�s��x��_�x�H��QV�(�8"iC�DC"�w<Gl�d��ۓ<5kb"��@�F
���N �LZr�ɶ��~b0x��J�8v�3E����!�۫�YY%/��0����P@b��F졐�'��L�Nu�RU48"���>��덐�s�R�2�\�vȹJ�Du a�� �s� ��\���5i�ö�v��<���N���HmpS����M��ƨ� "v� .[��E����Ⱥ��xi7�I>�ۇ� �:��mv����J���u��oqڀW�j���I`tP�i,Z ȿXSMqF��    IEND�B`�PK   <?XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   <?X��j�  '     jsons/user_defined.json�Mo�8�����)�S�|s�t�I���eQE%�ʒ��i��ޑ�4�Ht�nv����(�3�������kl�9�Y^�4�_l��U	7p�C#M��6�����gz��]�i������9<htk���NsSW�*ۺ*
[���B��:�L��9\�����!)F�c�4�	R	�)$��)��mL�o�]�O��s�3NS�E���1�)���DR��N��2ܖW0/�Iz�޽�B�]Y��m^��Y,۬�f[軣�h�X�P�#O���0Nvw�ԕ�M�'麭sX���j�>�Ӽ�����ței������`k
�����g�ǫ�a>�%c,�����{r~q�։�c���^�ƶN,c#/,٥���T�En�3��3�Ǌ���C�J���\P5�R/�;���P�s&q������_R7t,*�w���K����%wCǂ�~G)�б���)�)t}��M�P�Į�n섦�vy(�����+�0?�8\cm�u�N-�u��N����/t�hIOl�N�,�IUn�XcC���J7u�1J<���:��P|��,C'��"�(\ܓ��(]�V��]�'�-.6Q��'��ihc?��m^C�� ����5�&bW�"�G��%L%л'�ؤ�e�{[W[[���:��F�z蝇�l��v�D�����������=/����{Ľ��̛<)�����tC�C�o�kE]v�6mW�1�a�x��aL�J[���~��.n��}W�Oڙ�.��F�k;|ο��b^���6o���M׶U��Ќ��f���tm���e������-�D�� -=)�(2L"��IL�����-����85
얥(J!�.�6��Տ�ါ⡤��)c%B��#�Uw�C�"<g$��!��}ց�z�-�1S�'�:PGt��g����t8�]Op�Щ+)���	Z��^�{e�Nʴ��@�/"����d"��G�s�P��B&S��q��;-�f����^�ÿ���U[�K��� ׳Ӽ���M�����?���V�e]y0-�\P��gHE8C8�1%9�iL��N
����ĳ~+#m�ȈH,��GZ�BӘN�"�T��$	4�|N	��8�Z}7��鱇yx9u��/�J�/N�ۮ|i]Y����#�t�"-�A1Ilj�� ���O� PK
   <?X���A  F4                  cirkitFile.jsonPK
   <?X�����  �  /             n  images/37b7845a-1f46-4418-9ae8-cf8221840334.pngPK
   <?XeX�^Q3 P /             �2  images/a8051118-2cec-4f18-9b89-ac75f15be4ed.pngPK
   <?Xv����' dX /             (f images/afde01cf-9dc8-4de2-b588-5b54baed9cea.pngPK
   <?X$7h�!  �!  /             ]� images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   <?X@�G��  �  /             �� images/e086d210-4fa0-4a6d-a74c-91bedc336751.pngPK
   <?XP��/�  ǽ  /             �� images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   <?X��j�  '               y jsons/user_defined.jsonPK      �  �}   