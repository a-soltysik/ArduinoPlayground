PK   R�?X�O�:5  �.    cirkitFile.json՝�s"G�����Ut��m�31��ox�;�41jы��^G�h�%Z*�︽������\��7�?�7�����n7ۛѥ��w�������t1�������ލ.����_>���]���|̼(������zQ/�U9mǳ�b9�TV+��"����._��x����F�!���E�!���e�!���U�!���u�!���0CT!͛0CT!ͧa��B�ϲ������x��\?������b���2�i�9���Y�ܥ��j�������ϧu��YZ�'MU���^���E=^�6-��M����0�`;^�-^��Y$^��Y$^��Y$^��Y$^��Y$^��Y$^��Y$Z4� �����������}L�� ^����w�kx��a�L��a�L��a�L��a�L��a���0E�����9^w��"^;��"^;��8k��e�v�%2E�v�%2E�v�%2E�v�%2E�v�%2E�v�%Ҽ��ΰD���ΰD���ΰD���ΰD� ���kg��a�L��a�L��a�L��a�L��a�4��3,�)�3,�)�3,�)�3,�)�3,�)�_�⵳��ΰD���ΰD���ΰD���ΰD�O�3,�)�3,�)⵳'1�\x�?�a{K�����YmkFc_��_Y�(c}7��X:c�Ҽ`�+X�P:c�Ҽd�+Y�P:c�r�`��X�P:c������f�C錥�3ֻ	�Jg,]�7�w�Jg,]�OY怜w(��t.4$����E��,8�F_��_[p*GCg����Wt���ل'p:18��OX>���*Z�?8��|�����pNa��{xu(�_/DN�Y�˛}y��������g0�_l�G��`>�L��=,��|~�?��3�ϗ�g�������`��������0`��W��W��R����g0�/}�����g0�/ځ��ja����F�p�`���R�p�`���%^�p�`����i�p�`���eu�"p�`�����p�`��󥌰p�`���E���%^�5^p�(��Q����3���������3�ϗ�������3��������3�ϗI������3��x������3�ϗ���Up�`���E��p�`���v �p�`���F�p�`�����2z�	�?*8Tp�`����p�`����p�`���V#�p�`���&)�p�`����.�5�?X>���1��?X>������?X>�����?X>������?X>�����ԝ^���5�?X>������?X>���]��?X>������?X>���E���,��|����,��|ޖ��,�=�7�i�io¡=�b��vx�iԁ���.x�i�с��vx�i�ρ����x�ic͡�&:�㮷u���#��]���c��E��V���N�B#(�����kh	��>TC����OC���~KC���G��2����(�����{������#z����X�X�W�x]��_t�[;ne٬���MӯL_�u��go�I3��5㦘�q���xٮ��j��-�iUV��<����Sw��}�����;b����F�Q		%�$���AB���$���ABݾ�$���ABݞ�$����AB�~ܣ?�t������]�]�ge�K$W�����m�
7��� 1a�۰�M)�.�BLX�6��SJ��V�+�R�R;�}!�Ն&������LX���fCLX/�:N)�Ԇ��:^`u�R:l�1au���8�t؊b��x��qJ�M7Ǳ�x��qJ鰅7�ĝI�N�`u���8�t��b��x��qJ�8Ą�����a�p�	��V�)���V�+��SJ���!&�8wR��V�)��6�V�+��SJ�-�!&��WX��ۗC?�`u���8�t��b��x��qJ��9�������������a�t�	��5V�)����V�'X���CLX�`u��R�z��v\������a�_�`���8p��W�X�[�㪠��K.pU�WkvƁӥ�*諂��C;���q\�U��߽�q�t�8�
��`����8p��W}U��w}g8]j����*X�;�3�.A�UA_����N���`.P�����f����y��k"��6��c�eIoE�K��z[�󲤷��%�M�m�yY�[M��Ц��,�&�IhS�v^�%Hh�t2A�z[�C&h���6��}�eIo5qLB��{�󲤷�H&�M���yY�[M,��>��=/K����e���g��%���2	m��A�˒ފ~������,�&�IhS�z^��V��$����=/Kz��e����%���2	mz�=�&�IhMC��mOz��eZ�Ц�ޓ�jr���4��fWsa�&�IhMC�k�5�jr���4���Z�&�IhMC�k�5ފ�V]���e�&���\&�5����x��eZ��z����\&�5��J�x��eZ��z����\&�5����x��eZ��z���&�IhMC�D4�jr���4��E�&�IhMC�]4�jr���4�ޣF�h%�h)�&�U�\Vir���4��3H�&�IhMC뽏4�jr���4���I�&�IhMC뽨4�jr���4��SK�m��eZ��zo0���\&�5��8�x��eZ��z�6���\&�5����x��eZ��z�<���.�6�\VkrY��eZ��z/C���\&�5��d�x��eZ��zoI���\&�5��Ȕx;��2	�ih�ק�[M.�К��{�j���2	�=�v��g:���Q9�Mv�߈ʙ��U����r���@�3����� =P�L�硣���=���Pf���Zu�3��m`:T���.,Ce�A|n�СU�����*Ì�s�T�aF� ��0��܎�Ce>���M\��t���;��o]f��=�^��r�n���Jy�Tt2֎�EY6�j�l���YͳT�di�I3��5㦘�q���xٮ��j��-�iUV��Y��r�򩓙����bߎ.�����ݴw�����o�n �P�^+B	�nf�AB���"D�P�f�$���7B	�n&�AB�K$����AB�K+$�ɇ)�\���6V�+ܔR:<�	�݆oJ)�'Ä�o�
8����a�j�aE�RJ���0au���8��'&n��M��:^`u�RJ��%V���SJ�p&�a��x��qJ)�11LX/�:N)���/&�cu���8��}c0&�L
w*��%V�)%��1au���8���$0&���X���Ƅ��
�㔒��ǘ�:^au�R���wN�;)���
�㔒��Ř�:^au�R�u�V�+��SJ�N����5V�)%_��1au���8���0&��M��M���X��|�
Ƅ���㔒�����:>��8����cLX�`u����k�{k7h��%���IXM��
_{�6�&aM�ޚZ�U�j�4ﭣ�UA_�&a͹K�ko	= �$�y$�|q@�j�<G���[:�8�`5	k����Ӫ��
V���yo�<�
��`5	k����Ӫ��
V���5��`�I\Z�����oE�K�4��4��4�KBkZ��\�&}IhMC���k��$0	�ih�����&�5��a�x�IbZ���Z���4&�5��)�x�IdZ�������T&�5��������eZ���Z%���\&�5����x+�EL���&��\Vhr���4��N�&�IhMC�k�4�jr���4��&Q�&�IhMC�k+5�jr���4��FT�&�IhMC�k]5�jr���4��fWsa�&�IhMC�k�5�jr���4���Z�&�IhMC�k�5ފ�V]���e�&���\&�5����x��eZ��z����\&�5��J�x��eZ��z����\&�5����x��eZ��z���&�IhMC�D4�jr���4��E�&�IhMC�]4�jr���4�ޣF�h%�h)�&�U�\Vir���4��3H�&�IhMC뽏4�jr���4���I�&�IhMC뽨4�jr���4��SK�m��eZ��zo0���\&�5��8�x��eZ��z�6���\&�5����x��eZ��z�<���.�6�\VkrY��eZ��z/C���\&�5��d�x��eZ��zoI���\&�5��Ȕx;��2	�ih�ק�[M.�К��{�j���2	�=�v��g:���Q9�Mv���ʙ��U����r���@�3����� =P�L�硣���=���Pf���Zu�3��m`:T���	*Ì�s�q��j03���R9T�����*Ì�s;.�aF�}�~�2�����2���u{Ռ�U�s����v�,ʲYU�e��O�j���$K�N��լ7�4������v��V��l�N��Z=��,�c�O�?�ϯ����|��yt9�}��������U��on��ݪݍ._�������$f��xQ;]�w���}A�H!F`	����7��/bOo���O�O��o�H�+��ӐH�{���ſ�|[hN������XB�������u��oӷ|K��������D�g��a����R�ܘ�޾�m�k�o�3����I���,��?�L���	�#T�f^C��@�r 
`��x��1���>�����䞂-��I��o7�y�d������@_�$��7���0���3n}�i�S��=����A��	QЋ�t:̓����LI}ٝ�Zy���1�o���;�o	a8���p����D��쟟�ns�����vt����z}�����jt�kd��o �qa�����K��*� EX"uW�)����&H�H�U:A��D��	R�%Rw�P�",�����a��]�����Z�-b�O:Me�(Q\��j@y�k��e\Q��Pb��p!Y����ٸF:\�� *��6���E9)�����k�HŮ�X@��k��ՂQ��@��k����Q��@��k���Q��@��k��5�Q��@��k��U��
�^K���5��:�A� N ���i\�{[@=-�z��� POK���5�/���
��q��
p ���i\�{���V�+PO+���5�#���
��q�p ���i\���? ���i\���@=��z���X ��POk���5�G�����q�}p �t�Ӹ��T8�z:�i_#���Я��;4*99��"��Z7��{�u8=��`>��Ҽ�>��C�c��K�^�RN��3����Ŀ^_���e����ؿ^����e����ؿ^���e��K�^+QN��3�/�{�B9=�?��`���#��z�~���/�ŵ>nt�K�c'�FM��g��O%t,9]��
2��&��bi�pM�_�
2�	&|�����v%��CK8� [��-0�ф~Y8�!�]`B�	��v�C:���F�����l(0��hB_;@�ƦcLh4�/t�=�cLh4�/Ҡ=�O�P�cKAǖ��-0�ф�8����-0�ф������m&4��%��9&4��T��9&4�����9&4��as-�C:���F�"<�r:���F�B�C:���F��G�C:���F��M�C��/��/:��tN)�M�fi�M�}i�M��i�M苬i�M��i�M��a+:���F��|�C:���FzS�C:���FzC�C:���Fz3�C|�
�P��)�S*:���Fz�C:���Fz�C:���Fz��C:���Fz��C:���Fz��Ú�)0�ф������)0�фެ����)0�ф�h����)0�ф�$����)0�ф����_S�/��sJM甚�)0�ф�X����)0�ф�����)0�ф�Ќ���)0�фތ�pB���hBo$G{H���hBo�G{H��О"��c�!��mP���<�׈u�����5>x|�a���{�F�k:��^cϡ�'< �#��c�P����6T :
����q��F�C��㲿'�����=���q���vRC�����P�h��L��l÷����C� �㴿���]Կ��]��߶�fv5k�M1M㪭��]/Ƴ�j9[�Ӫ�V_{�gx�O���6+߻:����ϱqt�z��۩���[|����I����N��}����#�j�X��?����7?���n����#
?��#
?��#
?��#
?��#�[�6?�3ބ{�|�s\;: ;ww0�ݻ_�|g��}\��|����'٭Og�?�I�>�}���}��ߋ��լ>Qt촇P��n��>a��|3��q��ط?��׋e{���'c��������ò���w��*�w���*�wU�謁�-���G�ln�����v�=ˣI9/����k��jv�Oc�y9�n�{_~�������e��r�kw����v�ߴ]%����������~���w�x������w�ןݮ��ֻ�M����}�����Ϻ�������w޶�7���u��]�?w�]���>sg��/n�֋��ݮ�}��aG$����f�d����~��>��|��ӲyUg��o���}Y-�*�㦮Ӹ���x���x�,�-M�T���/����n;I�������� ��o΋�v��*����kovW���2�ū���1�����3�جxU��i����S�S�cG�L���9zP}t{ut{q����I�#�=����SMN_�o��'�ؗ{��1��ԦG��S�S��Y�����cztGst{}t{ut{q,���o�7�_�����f�e<��U�*�R�0��?f��t��8��a������g+�W��!�|��j�^5�Mg��/����>��b1����:>��������4īj�,����?k�y�A�m��n���>�U]=,��o�{m��#|�p:-�M������2JU�JӪ(Ӄ*Y�ZkRZ��TN�U~���ɲ���������{�|�YUr�����!�J�<z�SV�����f�}���<:Gee�i�Ũ��������>nV�w>����޵�{}9�Lӗ>=���W���w_�������7���Ο�[�C��&;|�ݽ]��)�?W�]�ɟ��n����o�'�N��Y=�"��n���5�U��a����ؿ�}�����s�X�w����[���������2����|u?�G\<�������h������~z3�������8��٠tO;��[�����D�G�&�p��k=I���{�ۿ^�ʦ��~K_y�q�n�w�e����I����&��;~T�<�W�~�j�g2�rqr�E5|��]0�:�����{[���9}���Q�e��{n����TA֟�n ��2�������9yؙ�P��Q����7���X�}�ow���|9����������Ĺ��n��o��������F��PK   �?X-Q�� �� /   images/2f436d2a-342e-4b79-b795-89e98e9450c4.png�uP\��7:@pw��������A��� !w�����܂��G��G���ݪ[�Φzv��տ%����E���*  @U��� �p  �L�WJ,�����I�� @��Ӡ��Y����
�

� ����r( �k����L  ��?���W2 ������A��E�zm���'�6(h ������UP��l�����
��A���o)��SPQ��d�`g��p�sr�srqPp�	rs��2A��K�?O���ի<l����U���Y�� 0����_�b^N@s[�le� By��NIac!B�ǣ®�$����qk��j��ؚXP��"	{	�؃݀^�v��^"��
�����()�bq���U[��L������"�e��I)�D!�ba)�)-��ב����� ���'�'������ ;'''�+����Ћ�������`Ws'7G�?c ���M���u����wRQ�'���?���6/�+;��=ۿ�pu��p�?�p��v�i�]�]��2`7���0��z'w��̱0gہ�_Y]_18�C��X��;���U���t�������g�/��/���-���/	J;���QOAZ��|AGs���� s^n^N^��7;М��������m	b��7(W7��9��+������A`n�9ȒӒ�Ӓ�ia	[�������kT��]�?P�P s�� �%����f�xyXxy@@�ς��/(sAYG{��v����lNVM�q�����%'+��(�v@7���9`�`�����)m{����?9��y�8��8�8��y�Ťvq}��?�%�_36�9�F �����;�\�@7GmGG;���?�U^�����_A�������L�C��w��������>��Y���U��_��sJ���������Bh��	�@��L�[������?�6��`���@nNNv>n?��%���� '//�%�?Q\-�<�.`	�W?���5*���?���?�=��;�����_N�d���l�n�0���3�[��S���Q�^+!�?K�?�����_!��_!��_!��_!������)������SI�� xyQ�����<l��dY�&�,;~�x��4)�b��M`�hd��R�Ϗ��,�,�Jx��-�������NNY���_�L� ��,�č�s	ڜG�g�͎?�ϼ}��y�@V�ws�?��9��zc��3�Ҫ�Yqlr��v3��bo�d��vz0����8�%�����g!9��wOͻ��?>�WL=�����T�M����Cm�b�*��gn-�$�5�m����NΎX�\�/}���eE4��b��6�@y�ھzѺ�յ����H��y��T�}x||�{1p+�*��_�yv��K?�)<�y�w�zN���jw�?`�� `n���fmV]��ȱ���D5}�?oF�o���������4kQT,�.{�[�[��z�T|iCq�7k��?և��䷿�žX�{��t���?=���X]B?x�c�bOķ`�t?/�<��C"E͑X�{�N�r��[���K���������z�q%$�t �t�tQ�\������UH5��T��; ;l���;i��F7=Cu�u�v_N�\�;�8#����@����]l�L?�
��%]���{�r|�<[z1J�[Bā��IˀB�����=l��xC�,�J���*כ�Z>��qKK��Hx�*�>`�.�L(�FJ��:W��JWsc����W��>y������0$��w*�ї�n�n����_��W�L����ʘK��щ��=�eZ��l�9L�S+��^��D���Pm��p�N���WP� ��cNK}�/ļ6K��o�Įo�=/>��ëݶ\�{���V5hڊǲ��&Ӏ�Ό�
����A��z&��ǫ�c�7 ɋf�=�|W�F��OS��'� ��Ql���;�Nl��K���}2@�Jp�R���ʇ��x�Ǩ��f��W���I�oC7?ɩ7�`㛤I;�&R@��8�%��j�������9[@��r!&ѷg�,p�~�at�U�;�E����g�i��c��#U��������_g�O=/�����%�֊�g�[��[����=�6v�>��_9����ŰXM�`y�@��=���'������G) ��1��)�C0�P�L� `�����8��z��P�e��Ę�9!���Y���^z)��3:����^��e"��9��~�*�����81#lt���3�}-���zǌ���xI颌�F* Ej"`��{8J��s����|8[�����ǌ���kx�y�axd{�[}4l�kx�맖��ΗV)�v�[i���d��K{W���0����1��莉�%��19���F�����0��0����n���&d��p��j~t��l'/{� ��I1'�4�QZ+(<(�J��7Z鵪Y'��N�pUQ�@ͩ7�*�������.��<����^#ϙ�.vH�	�5�� #��w�-"M�G��QI[ ����Ϫ��}�$/u�m�ܯ�Ks���9���4�fݞE�!��]�es'�CGOB�i�Ò�jg'/9m��/g�-6�/��5˨'J�� �ƮԶǃ��v�1ߕ���k��R<r���x���݀[߀՛������"t������J��|�S͉���(J�j������臇yⳎ�\�9(��5��2���KQ#D �ϥi�=/��©��
{'�3�%J��DOß�4�'���Ёļ[�EIHOА��3�׋�	B!�Sb���PZ���v������i�K��st4"����k~�B�@�� �܎�5�����7�%��#'�F!vccME��&A��y�zYW{L6��k�Y2}�	<i��y>����{�u?l��nj�7Ԯ����=����)�谕T|��\�Z�9��D��W�V�<#�PH�FW����M�C��a݃#k���ْ�Ҵg2 �=y�꥞�������.��q{3�̜�>���Q�9��=���t�`�}jl7\a�C�_���g"w(E$F8Z���ٰڦx�Jþ�� �S�E]PQ��81{��D�$Smk!;z,�����4RR�C���w�*(D��*.�4,�x쉂�;_�M0�Ŏ�Y\��2�o��=Mq����x�˹�=�y�o�ZĚ�c�M�`�k�yX�}vK�|y�k��i|�����.&���R�<x%����*f�̈iZh%��6�,O����̙#��} ������̓^RMM�Ь#ۜGDHdsS\xf��,ֆ�}��&���.f��>�����=�]"�KC�R�ۀ~��B�K`�u�m�~h�,\���\>U@��0+Y4E�*�L���4�qVL@q�~k�G�Ň�p�[R
uf%��բ)�an���P��/�v�p�t��_B�6����	v@@�R�i঻��}Z���][�����ˊ\���c���u���Z7�
�{ؤ��s���i��	��G8j�ï��+�����U(f���;C�l\D�kio��5���+w`0T�>A9)#"u���D L}�B�!\�8��\n�d|ŧ �uI�P]�������c$�D�¨)�`L�S[��~(lL��B??�/�{y��@-#�w!�l��5�?��!v@���@:}��O�/o�Ḱ��o(b.LP��V��j��z��$v�3�W[_s��&�?5=�?\��x�p}i1-�c64�0��P��eы>�L�^Y�J��}�#����:�h�I @�Eo�xU��]�~�Q�;�{*4+��"���3�(&'��� =��z�L� �@|��C��v}�E�
.�'OA�6�O��5�T*�/��7�lx�
T� *s>���K�)���ݴ���iU@��cwٚ�I�0�B�F�|�2(�P✳r�g�;n?н���&RV;��"�HV�s�V��L��D�p��j��؞���:��Oo4��l�[L�/���	
6������f�Xi�H� �\�i��;�
�q �t�����j�nq%�D�[��Lw*ΉA�b�-ĒC!(c�8
f=����?��m�WO�*�C7ʗ��Z�>Xqm����i'���?��������W� ��������Mo�{n}��3�r�q���LĻ&j��,��BWI���+�xw]��BO��x>�nfa�,έ�aV��s;�a(:e=�7���zzz�X�j	5���^�H��\oІ�4�xM��~c��hX�~�9�	�kߴ��r<::
f��">{����}�<��Fo�؉����K�介���#�r`D�؝�L�	�x��J�^-5�����_��M�d��k��b�,G�nc6�	����Um���d~�ǆ��K��9A�"x�&��L	����,v׮�B��NO���2� �>hpE8��6��l�hz/��{�e�5X/U>�K���@�2e�d���\���|�����Շ[WD�����:�n�ǓQ¨�FC�� �TgȟAU +���e��H�U��
��ˏ��̬}}j�nts�WZ�N�W}	�)�e�e���;r���Į���^�_*�p[�~�B��<]��wr��"'vO���H�c[PD_m�=�C��Ø�q����8uQS�W����^O�[�'4��L��@�����o-� ���2����'UȂ$k�Ga0n纃���&�,撷����"�h�5��em\ ]$ݚ�.����!�aR]vo���z$��4�V�Uσ3�����A��%L.�N13Y5�i��PP3�3$�3���UG�̙�� h��y������]#ː��7�}�S�?��tn�B����S�SV�&�ҡs���j>��=$f����-�Q��E���W�����\LP�>��i�a۸��f�����e�4�Ŗ�v!��W�W�6�l*�� ���Q�lnfvv�ңp��9�,u�F�R�_�Ae���B��x��Jz�׼#s@q�7z������xs��4�h�?%0d0?e��(%eI�!�I�m��p��7�&7�[��33�5�el�-�~��b��@�i��S��2VU�C�v�č��.����!\=_e��LD�3�� �5�I�P4��*��������Y��.���)�@�L6���!�#�� ����Չ�Q��C"�/G17{ϳ��'�������q�oz�n�/��aK�(�P੽�#����e��c�Xr����{]�'_ �	)2>S�z&g���`��Ƽ4��*e�;�y�Q��ޡ]�8�<E�0GS�EFA�]'@.��-+k@�����EVH��ەg`�-��"(�'���R
��ڄ��M�Q�m�H�ȭ�{����ǋp�D�`�F�*+�������H@��։��Z���6�*�D�e�>�v�ɴ/x�g�2���2
��% go �	Ɉt�֊��a�/Q�b�kxI8�+.f�����.�T�)|�.���x���go��uKOч��痧=�����28�S�x��3	1͠s��K�A��	45����07����@�<�k9q�tM�:@�\]�;�g#����g4L*�=���|S6�c�u/�`��"HB�Cq1��q̡(������ߣ�Y��Ȓ���ҷ�~���xZӈ�R��R�6��-����3K.z����:����M~s]��õj��ޯ?P:u����h�muy�فp������ێ$'_�
�s��:߰�jAT��inyIg��i�۞������>C���=�tt� .,l���sXqZQ}���\�P�����;���aGQW�~+��w��
�3���\$I�/��%�d*�8��s�R��T���|�٧U=��;�V&Es��՚�?g��Usw��]��T��p�]r&���:��y���4@�)���aҼL�t���g'���Fa��p��6FO��]�<�LR�Y��5���`�耜,�tC�>�������ߦH'Й���R+y���� p���K��c�υ�c�R����-������t,�H����f����}����<܋�L��54z�k���-�U��xp"^�)dҴ����zP�PcD�FQ��ZP^<9K	V^���^����"&��8�5��U[���AJ�2�~��$��R7xR��q���՝FJ�꣮Ŀ��W�̳ܠ<l|�t�������"�A 	��O欕9FM|>��;���;�uϓ!��p���д��#����J�/
=F�(4_Ԯ������Z��u��SC�����%k��b@(O@��f��R7��D��(��j?X�;����&����`����)������7ϔio�40�Ho���7d�z�aq���\d6�W�@X��2����Ω�;�ӵ!Pĩ�#�Gψ��0!���qߝYj�I*������-��J�ߗ��dB��+"$�?��}����d�)ˌ)6F2ޏy�8��<�h���t��i#��;`U�D����-��2���ߨ�D\���e�J�[�xzXg��	� ;<�c����	�D�c~� ��}��� =��ޗ�t������	_�����>!����:�c��Tז�	�.�>Jj0k�KN$�'���Z��Z��֤������DbH+�$f>�ݿj�7b-��T��9+�a��tFu{�:I�4w��tþ�d�<��*/�<������N���棃:/`�!R��ST/�73GJ�'��C��U�����B��֡�F@Z"#Ҏ:�/�AJ����SO�s�	`{�U��2��[�0�E�,''�,������55xuj��~7`�3��506b_*.Ys��(��Y��^�J�z��#
f�"� 6��IG0@_���JCel��%� ����2ɕ�R�O���zM.b l6��ٚG�_~FT�����	�GoL��ں���(�F��b�q�/��f&z��0ڧ�p^&vj�d��`o�<��&*�΁ �+[���m<SX:��k��u�TΆ��v�}�}9�U2�Xc=�=3͆G^�& n�z�:*��;��Q��a���IvL�􏻽{�*�9���~�����q���+�֞�^0w+�i�*�,�q3�|0��m��x+-��CWHL\��t�v�Ʊ~��*��y���X�E#��B�K_<��E����A���+mh�{ܗ���&%��׎����g0�rb�ۼ�!��"�4�q��u��6����� ����<^��!�{���	W����>�ޙ=���z�vZ���aIpi̊U�K\@�L)y�R�ɄW-�=���*L,fS�2`�z������SK<�`��X�Hi	t�gn c�~��L.>����.]Ի+�޳JN��������U��3ǫk8s�,PW�����mM'��'��Tiw)w ��@�~_Nv�4[�-�9�~E������|4���2嶫�3���#�r���+��'%�Z�
1��ۅF9`ٚ��l�Ω_o|Ҥ��|��C�L����;.��A��!�Ed��\�@�]�ۖOs��X�GG����X�����1k��I�+Y�'�&Y��0�Zb�*�k�9�24G~=��8bx�/~_P��8h�3��>?���V:-A�&����Ͱ�0�g�C�7�- Ɂɼi����I	^�v���_d�.��<��	�GGm2	� 7{�]7�~*��(� ����`��*9	��Who���'/�(����iv�b������?���b:�w��x%��� \�DӺН���.sI�#�����w��)��M�@p@.�^��\�'�����A����Pʯc�F/4j��'����2���!]nV?���z�����X�Ǚ�h$HU�/'r9�v59�˭�t��h*�<�n��'�u���yd�-t�h(������ωBhE3Q�ћޱ����|SiQ4����̒<��{Il2�b�s-:d ��E��^YF�3�]�O����6��%!�/ǥ P�L>�P�D*��#�1d��7�0T1۰�f]���|��E��/�^-��� R#�j7�8,1Ҥ=�z����;�\P��e6����$`�sb��v����Q}�Mi�9�zh<!_`�g;4~�-ԏ�r� Ϋγa�Z�_��%�i���S��0�Id�T����OnN�����7꼳!ZP��6������H� A <���yg1�K����x�{H&ޡ'�p߇�ҭ�+xfS3�b~S;N�V�9W��=����G�Z�,��]�F�Vm�ʦ�~U8�i�mM0X7�UrCɴ�e�V~�#��Ҷg���,FW8����`T�u\��>��J)�����Ɓ)����!^Q5�#8H��k~��%Op&c��DDH��
��0	�o���		����Ր�XE�������Ү������`n��S��^L-g��o����x�����!�P^v�#Y�A֣ӗ���|Ͽ)��*5��w�p�G��B�-��V� h�<�\��"�`0��+���i>��P6������5ǌ�<S��qa"��I6���@�j2pC��ν�׵_p6�q��f���P�E'�"Ͱ��� ���6~�g7`�K�=�<��&E�<�@�ڝ�>7��"��3z��:
��^�r�ntuɐ�.���V�eR�"���ONNj�	2�}m"��WL�T���Rd9�;����FOڟ�On7��o�NC���#� �p~�Mpt��A�ۦ.������>�����F+��eI:\9*��&�w�[�2$��wl^�@y��sͧ+��� bʣ�M濏)��,8QC���Cov�8r�1ͪ�Q��/��]�(7�����	`��t���!ua8wNx�Rj�~�
�6�ؙ}�E��osi�'��A��A���
ڸҙ}�e�%�#���������Ne���'�#�����EQ�$����6�Vϒ	0�	M��g�l��D�Ņ��u�!,L@I�\9�i��։.���`|�W��TJ�*=0{���uCi�����)ܶ�*�\��Vp�}����:ԁ$P���~/�s���0^m,a��%�\AJV���<�]���6�V���:��|[�K�k�3�+����Z�^�m,Lc@K �?ǅŁ �&#	~�����~&5Ǟ�bm��t�-�״�z�e��s�I��&	��EU?���E�4��/���Ex�/�����K�3���H�T�lw�h��:�����4|*�<	��P�2���O�������O�w�י�5��)���X���V�zI4��ތNY�������2gW|��ś�9�ojX�)�,5����+d��[.|��y?1���-2�e? F}�C��� �}��'���4�C���8����+(������nu��}%�Cv�dTj,Dŀ���/�w�9p��E�4�6u6����=F��}t8[@�Q�B�m\?�zҿ�Nﭦ��Ǹ�M�w��R
�L�#�\��f>�_�=)<���}>87�ߒ�J>|��h�"��C��?#��K!u�+��>5�%���4#I&�}�M*��^N�
�(�F���Z6�T>8�}�!S�'�cR�$�.�1������s����g^Ce��԰3
��f�-��h�D�xgw�n���<���!��Suk!0�{	=\��WM׹���GY�NB��Ŏ;q�jNRǰ|�"�M X����#��g�ϢZv�h��\��;ݐ��2��o=�C���X{����WN�}�H���������6�{�ȧD拎s��R�u�Aĉ����s���i�'=�J�����v���6���+��L~�j�8G�9�;��r�[C�a�NI,���|B�D�xw��"��m��F�(���vQi��)�C��������9�G�"ݰ�׺�	�!в� *�D���.�E��H�v�r�.Zl"�D��'�Ƭl9���lP��u�Y;�l��sVؐ�U�M�D�pX逊��?����SV.�ذ�I�@x��.s6=^}���8�a$�t���J��Ma���xy>M^��Y�;�&��S�u�,�_�.�!Q/j��Tz�JY�@�?EB-8iہ2�kǺ������	X$�$���B>���/u*����a��@4`��	:�i/�B���9~}�R麘!Q���@n+L�~	o{۴]�����P�6��OSIFf+����;q�.�EД�6����7� �2�Ѻ1��Ti���w'��O����h=�Q'�)���{��",eBW�.g�����щ#�g��'?��Q�e�����E�Pa(*y����9��Yd��H�r�Ú������A�k������i��EW���<=�II\�m����懟	tTZ�����Fی+��-����"�<�5#n����΄φ��\�R���N)`.��_=�GD�LY � Y?�F�.�R�8,�ܺ�b�����
��|/�7�b�F�s����NR�)7:�0y�	sD��P�D91�L+:k�bX=/n�њ�D������^����ĸ��\#a��^�^��^�݂�q��(�<�>���� �T�[�L�P3@���ЙA�oLF�h|pN���X������G/�Y�D�u�Mt4}C��{ۓo�RU}�qX����!r�G�{˪&�y�t{���5?�7��fR���e��N�f@K\u��=y��{��؀�&�%� �f_���
�G�k&����D?�w(��>��e�GD5M��kf�V��"��UdE�Bn�Ba0��	9�[!ό*L��N�<6[��e���w����h�%��2î�v_~�;uQ�QÝ�x��6��R�{^�'K�J��Q�y��E;�ŏ��8�߉>�jW�nW�����Qˣ��V���ޑ�=��,��r�}*�})�y�����ċ�� �̩3���T�����(I1Ѐ�Z��,�\밙y1SG`��K���?X[A��O����~f0������c�� T����v_�
G+/G��� tyK1=�I��s����ZC��%9����
~��G�I�*��8�!����u�fA������1S�a�i�t���ᠯ�!��5u�j.v̙�W�Z}oL�d�ߎe���]����<��գ�:v�d��!������c���M���^h?�����rg���ĩ��]��*��/���!�ʌ̥`du!�P��y�8d{�W���K�f?�/tC����9>[6���@<�����Q�4�f��~94�H�i�X���6���t�d�#�]�B���W�+s���!�F��]_�<�!�׭��,���O;u��b�Q��3*o��֔XD�a�J/����\�(U}�i�`�S�(H��z�d�0i�t
]�|�[�2	Z>7�d���k�<��AE���?��"�!�>� ����8������}�����oP�fQ�����X���bb������U�xr��Yϑ�>/:l�}np=���JOg��Ϳ)�l�K�aߘ�&����J������*ZB�Lj�y��ه���7�zG����`�t9Վ�D�R�rˏ"��A��r��<���}a(��	4&.L̈�X<y�a��/e��A�8�p�uiɰw"�)�mW����	Z;0N�	�M(����� ��Wdi����stg.�Q�g9@�ƚ.���=O��.<_z�1�q�_bF#��T�@�|86(2�h��n������ �Tz�5H�z8X}ώI1��f��`ߒT͐Z����+t��3�5�u��L�h��M�M�A;	��쩑���'x��o�4Uy�:��-#<�\�;Ld-y���#k ����o��p}�u�SP����J'��xJ�����	fqu)L턾V>��tJ�{��]�:��һ*͌AB8�����m��ɭ^�V��k�e
3G�Ó�8������h�d�x�:�UIl3��� � �L]�[@{?(��O�G�c�*��o��G�xǒq�U��9��7M;�F��2��/ļ��LfXޜ�<�f��6�]�݃]���gDզ�	���_��mdj>��-�΅-�KQ�u����6�6�Η��I�RgI�]yS|!��;����bOW� �`�K���
�����ϊכ�`�x_n�B\���q��u�S[�Ȕr��H����u���ht���D�)�b��"�w֪eke)� ���JM�	Dn�}��*dz�o���'�!�=��U�����<�h��i6>n1%G㿥��ّ
�Ea�fA.+������ߋ�->����0�"8K���"��ShHN������0;q]t�.�{�3 *,��%`b��㻎BӢ�'P�}VS��ۻE$%-�L�*�z��-O1��6ϸA�s����=]YQ��o\Y�]�f'ذm�(i�f�k�'>��̅SU̓��vYV��57�mK�d�a�놝K����+���D�ǖ�)�BR�2����f}�VIg_��L/�����G���F��N�F:-�d�ۘ}���oڍԨ<vU���m�f0VX����v+l c\�؁(Y�6;`יV9���\�n�ؽ�=&K:|+m�]�$)K,�I�������SEwx4#G��?�K6���/�-�1�)X"�W��*�+|����*���dƋ�mLf���W�qO'�x�V3�t�/
	;'���:�y��7z �|l^ˏ$	�N�Čdy[��g�,'�+	���L)�ʹ�f��4�E4��F�*�*t�����(�	�5�X��?�+��V5�´E��x�8�K�vXr�5�z��$�m
��O�Rع�W#Q�����}u�A��ɒ�W�wt�C��n�B;s��&	G3[���O�s�m���@�G�p����:�z6�Y"�j�W=#����]k0ONI_`�P�ڿ��\)\`�e�@�[?�xqJ6W�X��e�OXZ��例�ɖ�5�����n3���w^�˳S��%X��T�I�"|N�\l�SL����w�7�=����*�qZ�^��p��Ӳ��^�/C���@�a��n�޻�P���}ߖ=\�
{�2����]>�6��&Z1��ꪮ~���sb�����2���G��0Ԭ�ԗ�`��(s���%ج�
��t����aT\���"�Qޗ��$ZOBe)�Ow�BQ�@���X��SŴ�h� Z�T���O�Kj���ʻM&�EB�=N����^�S�@V��@���z�bM~�W�?1�}"� JI\N�	�^gb��DT!�2�v��6�B	���.U{�=�a��cV�~*���$�|��%:�X�H�
�՗ѽ�1
/+�Z̠W����t��'c�#�FD7y�#�Ȋ�(c볢�݌;�L7���q��@�W$k4��U42���B���֑\�/d�]_e&��vN~�?S5-D��=3C3���W�QVN�������F���Q��ЬK�$:�~nF�v�5��$�Tji����k ��-�yh�@V��?#.��f�Q�k�0;o6�.]P�W$�Η���	�}��|V���6ߡ��,j�C�7>�Ya-�,S:C�A��־���mH<T0�6D���w�~��t`ApD�^�rG^�H�����(�b�v�se��!�l!���'��w�GQ���<T�*�D���ן=N.*t5z=�p��qy&<���^�7�6�=�DOf`8��[�f�a�H�.Q�4����CT&/T
f#R��%�S�B�Ke6'�*z#+<�Ү�FXR4�#$`�� g��%�e�R��V�"V~�d��Ce���9�)	�i5W�.V<3���^�c�o�&��M%Q9��2�o�_>	�������X](���;��|�|l��3f����6�Xb}@�����p�mj��4�Z�>���׊����Z��]�^tGf�z���t��t-+�i�F���iO#�t�|*зg�%�UO�&X8�/�M���n��_�h�6?=���ތ����t�YYv���t�d1��U��!���"J��,#�=�7�?�ټ���+�Sqg�U��$2�y��]�&�8:�4�R�n�'�:}?������G��гC�L.�q�Ϊ��3 �8�=�P��T��`嶸ǜ;�]���s�Gb�s�/b���1�u=�z�6��N1�"��c��z�b/c���Ƥ�"�H��_��N"p�x)6tPo�6��Hf6�v��m)�/f��뿯�5'[���zܜf�UU<rD����N9��d_F����䡭�9���1Q��e�`Z�U���L�W��E���l�K�Q\%��ĕ���h'`�i5�p?�Q���F~1`|E���8��:t?h��bO�<�f�|
�����U��R���T��f��lX{Ϥ��[&d
��i��g֚uqj���e�N|�vN^]��o�Tc���}��][�C�j8Q R� �R�<5�D�:3|Y���9�ҧ��f��@���&D�*>O�;�B��$���1��K�8��S+�Cxn+s*m��~obG��f�;��m��|qK�酔o��ժ{mK�aS3S�gk5[�O^���B��u�׻HfXU�n����ϴ�2r2?��BN%���š����W��8�cs�d#F��1���3Kl7,>���PR�Iw���]l�ᚵ���[3����X�8���2��@���� �9�G�E�S��kV�e���Ը��#��w��1�N�G��$,�]Q�p����2��:F�Ka�Q�\��{�E���r�]--{�ظ*6�,��A�s|d[)�0?�5�0uy���}��b�z�}`4�I���� �<���*����A_���/���{����T��l�����wX�d쿫fF�κk���1�B%:�-h��һi�љ���!�v�i�J�A�L[E؈r����o*ĴЋT��.�ᱣ=�u�����=Y�c�rU;C"hzIߞ��+i�q�.�
$�k��#䚚W):�>[�t��/$�^$��4`�E��G�c_��i����I������.����X�l�h�'>�
q78�p(G�r8��,���C�|fU����y�0ߡb��v!����<��z���y�IP0�ɝ�RA���pۥ��)�*/7�=�@a��gw���m��{K�_M��٢AU��`C_�y+W��<9�Fq�0�lRƌ s�YiE_�k�D٠�]wyt4��ݲ0S5\No]
�Q���P7#�e��DMI%�N��X�8D���f��gN�$gכf�g���*���*���+j��"��-���bh	�PtW��'Kw"~�_X]��:��S}/^�0 �ќ8Oj�b��]����`�D��1��-p��6ra�撾W����L3��1v�����O6�M�.Z����,P�p;�޼(�6�s=��2wƑ��Fgf��K�E����f3��mzz�2�R�����4D�o�D]F>�Ӥ.�Qz��������3;i���ᔋ�� ����:o�>]��~��;P����{�v�3�nHa}�/bU��$�b@��'��<��T��]�68�C<�e��H��\�����������;��A����3��ö�y��Jv2e����!�m�ܣƻ{O���r�ݷ �錾�vD�������$��c�:��9E�@ݾ;9�t۝ҴL�N��vH\�U���15��GȓN"1��6A-�kfu�J������g�OB�QT��H�<��y/).��.��ٌ�+\���xH���m�W�m����`��'y+��eiAֿ�s#�Ut�`���.o����i�S]����Z�\�t���T:J��kx**�B�/�z��H�������in���f���FiL�rG#U�Sn/���!^Ƞf�Z:����������a(�[=�]]&s�Ο�Q;"���C�uU��u��(� x��$����1�{i ZLHרblu&i�{�qADG�[�Ō֘���]�6���|4�+��,���
/�ӷn�c�tU��_��x�&L��(E3?f�8�ǒ>�_��lB�P�!]���1�-E�KeJ�S�9ki�.߅�(�B��')n�s}W��Ol�,��Qɟ�IG1S�7��l�A�Wºo8�򕂵G�h�Ȱ�[���9;��t��y�)�����b�ǂp��Hc�@���aÖC癮����(�e�7�q@�hL���hq�a"���;�Lu��tŉ��xu��\���EG���_;��r.V�2u��V�ǉo�4<��bj=G6GT���}�ӫ�X��5Lg"�[V]P�[�7����Y���Hc�0?�~�W�^0�ue-����2+(-K*�$Ah�i���xT{c'�ŀb&
g�(^�0�)�s�26.��:מ:2� א�42	gI��>��~�P�׮X4����W��br��-�p_^��
sowG�iG�֌�#˂xF��H���:��Bm�(/�V�Un7m���X�%b�����ˎ�{���-M:��G	"���'��
y����h	ru^��ص�f ~�Ɂ6BM�L��gc��.��۝*��*S1��@,d%Z��6�n�_�7"�*�������p�|�rݱ1��c�]�~	�\x�)�]�r��kl(r�r�'�GGP�/ -@ҿ���Ԝ$�9fc��{T :�l�\���m��iɠ�i�l�.'&l1I��Ǡ��z�$��1�g�\��j� ۛ�z�\c��8I�d��@\2Q@D*���{��j��V:�P�zӖ�u�]� j��� �)�6��&Ӧ
(Y2�ʿT��ik� .�ٞN�\xbY�d=8b�;{�qNdB�1��v�֭;�Y����Ϗ��������9�� �L&������P���﹜(·}�J��9��XQ1�@�\�8�Aj�y��b@��@�K�w�����צZR����p�v����.��k]��m�P^��<�)��X_�;�7�Ri%M�l>)<=�%�g�,���\�OV�Ȑ?f��|2��΂^�٣���������k����lr���j '�I@�3�9��g�a��B���2>g `�
|V��/l�_�H�{���,3}�gs(��T��e�:��jp`[qS��*��bT��;��5�Y���"��-�<w��G��Uguz����2yT!K�UZ��'%��pi�ZQ��p��f:�A��"�h8�=�9��v���}��A"Y�E�AZFJ�����5���E�J���fCS&������ޯ�iX���-<l%���3�Ȥ�uK�ɸK[`V>��*�d7�L��{�Cy!��iޫ��SXd�_�/^�2(TJ}q
*|Ngf�>����8����,L��m���u��a��.Oh�6L_�\��,5��L��^ ���H�#���rO���93� 1�u�����.gb�v��m�*2��J;�C�%o&��"Nn���i�b��2�S���q^ŇJ��'t�D���~Ʊ�����
�Oj8t��إ��}.��X �҂��¾]d��'�4��s�w�l�Am�)%Qx̲�!byo�����>9I59(}�y�>%�{A�sY��.X�"�
.� �u9�~)�	S�A����`���+��?�k�<7��@bJ�J+�p(�?-���R�Ս@r��,�( x�v��R?�"Ȉǫ/��h8W���I�4	R�ɥE�a) e�眳�������[f�Ϧ\����=�w�Uz��1=y�����ǂB`8Oɥ5�dx���p��dȟ/���{?+r1���h�-�1h�1
��%��ǀQ��dP�wxxHGG�� �S>�L9���z�A�� �Nu����9��@� �S�~v��P^� [5W��?�6���M&"��
�A�Vi&��ռ��P�l9�@?'����k��P�������Yl�@g1\ɫ��Wb����j����|�=p'�q�Fþ��s�R�{8@��+�#�'��G����Gtrr�ޱ��os�����R��3���Jc����aN����_{I�MOW�d *�����6P@��0��S�����-H �Yg�Ԍ9XbP���\o%M9S�z�a؟�[ݠ?
��@pq1�������} pފr�~$�(F#�3��(���a0ᏎNX������Q���Qh�T�р9�+��W�@�����1�.D�M� JfV��^
�w�$/xb�n}EP�h���I߷:�&m�Ԏm+�81G���A O��Xt��Փp�_ ��(���Gc(1{�X�YLAF�1�<���p�0�å�ʘ��!�������օ@9��r]�� =���c.��4��5�F���ͦO�˘͖z?S�ੋ���"�H�P��� �c�P��E,�(�{j͢�s�J��.H�&��3��a����ܴ���/�H�(�k.c�<�c@��~Oc{���o��@L�!�Z LPp��9�;�̡L�gtr|�j^7���)�`���i:���,8�8  �\$LL��9�%����〘rttDx������ko�o����(�ʽW��\�t����(�ېu#�ٔ��c�|���6%"�������(��/��w���8��r�2��4�N %�8i�rF���@¡4t ���Ym$�t#�,��p)6P�9�q` ��	�K���g*-��@�LY-h���R���ͷފJ�2��RJVR�g8 ��lN��G�������<x@{����g��u����m���wigwę��<y�
�W� ,�N�@�Ϧi��z�T���*��90��K�k8�.K�ۡ4���oeI-�;mC��]˟��=�z�e�6�P:h%���/�k@Ճ�R��{Q���Z;�I����e%)�c����{/��`�}\ (E����k��:Xx?yB��r�^}�����l4��h���U�"�tvw��E *��XB�$d���R�����A+�ݥ�w���uD�I�3q�y��Ɯ�	�vg3	<\,�f����}0�����_��y�e�й昵Ԑ�9l�f��O�]�Iu?S�m�^�Ģ���B�V1G��f`�3��p�-�.�u���c�\@ �Bt�����ŔW��p��xph��ȉ��+w�=�yM/Ni��t��A �a��sv�'�e��2 ����:@@29?Ǟ�2 6 �r���]L��>�õ+Ρr�u~��$Xwfl��T��@�0����oS�����m��;iIf6���F�Zퟁ�\��,B{h$��8�+B����5uA���'���&�M�P+ypX��
���d�,�0ƊcX�pX�%Z7c�e�	N/��p�$�frq���L@ir~��cpd���4�}D����o��g���ׂ�rB�� c����Oyp^L�Y����X � wJ ��ï�s<�Y p(���_a��Xpp��&|�/����WY�rtt�<	�u�z�'�3:=;
�2}U�X!$B�
�=̈́k�Jy�S�q2�5%�Q��T�3�,o^��L��>x�18����	�����hR�N����X�v��kz�$^�ƞ��V�K%�cR�顚0���l�+�4�9�i�h� %.��eA�x�%c1��I	]D��T�4 ǲ%+0y� ��"D��*5ON������D�j���E�X�3� ?d�gzqL��	��<$�	)�WOr˼&��=z�@S��Ǚ@;9~��H�0�%�����k�	���M��׿T?-���4��0��+�ٕ�n��xqk�IP�	���ơ�Z���"Ы\I�o��$YJ�4Sۯ$M�(�\��C�,,,Q�f�R03��L=��9e���
L�aˍCKR�f�vh�g<��17P�$��ud���,Y����W���f$y�P87I�uk��N�����BĈ��	x��H% �����<��$x���\���.�jx�Z鄯��
{M��i2d�%�Ɖ�4�Tn��h�O&��t5����&{Ƽ�T-�x�嚽��T@��2�4�~������RX8^��%{�BW�:�V�"�E���G5)� ��� Au�`Nz���<|G��A�3�N�DܸIGU���I�h��q�+��r��mE�Ds�T��v���qﲩ�V9�vcr57��z���U�)L�tͷ0��M}q&��\�/�W)�F� �`�0�ǱToR�>%�%�pr���pngn�&��`�J��A1�"�Jr( V$yn��T�B����-m4,�q�#��V����g~1%�8UV��ϣ��M��^j'5�C�ۅ]�۱7��U��P]��E��ojFO����V�'�N�y�}\�M��(�gc�'��6�
��_��������X�t6ی'W�z�e �D����Bk�I}%h!�pV�q��:rg/��-3�r'�'gI��L~֋TK��	6�]�jj=M�
F+��֫ۡ�>�J/!��DL�CSKa
>F��E^޻@[ǶL.٢�L�~�SI��fO+��+זR���A��ZfԳ���8��7�81�U�ɐ��D��:n�����U�P3{��F�¡�� �����ԛ��Џ�Y `���|'2ֿTlj��
��^�t�zt�K�w_�v�r))�Ҁ�����e'�l�r�l@Y!	,�\>�:�P�R�!���z@�g4ȸ1��Y'ѫ�<L3�>�8n�r�+�)[�������vG ����J<�gA��Z����i�@c��ixѻ���/�t^��C]
ش~���7z��s�6Pa���[��ī�r�%f���쬌�Od�h��R��:��>���[V�/�0�(�c�5,.��Hud	�$\��sv�+Ey�ܔ&��4��0 Q]���`�rm]H4�^���:�Tq��n��^ѯ� %[�a�Mں޿S�U��U9�&~U�I��������_�W%�[(_�"�s���@��q�vO���q,�8exw-��k{U�2סK�(�P�JZ��I�l$��"�g�������6�?e�,�����Q1kO�堎��v���M9��v�ְ��`��X:�M���`�F2_%|U��C8����oI�$�05�1��t�,X��NFѡm�h��q�W�ݾ����6_��j����8��R��~^<���JW����q���
����p(Y͡��F�l$�)�z����6h��E���+a.?�D���[+U���ă
��\���%�.%!�N�*zU��?L4"kn�9�S-AN�'y�ΌT�,a8&��5�ަ�iN��an&#���+ ���r/�7:����8����ŏ�:�K��E�IuH��@*j��H08O�vT��o=����d"3�h�uԸ�JV$�:>#�!Wǡ�LX��$��ӎ����?Y�����U@�n�^�J"�e�kɶ�*��m��?�AY��p������ڷW��k|��ל��t(�ӥ����z+�q7�Y���s�c�˲
\�6P��2�)�x���\�M��)x������u �	l��T��A���բ�T T Q��D9Sӷ��LW�X?�G���R�R�L?� �+Yt8����t�� ǲ��m/�xL`��"-@�o��D1������������</�D�z	�⓯?Y��hq�㢖^S�;���e]-��x��0�T%��$�]drͶA��1��d�upc�e����+�ae5P��k�8$�.}Z���wb����ۡg�p�i(ϝ"K�Tg:3��^'�T)\����}L�p)f.���wg"�L|�d��VK�=���d�H��e(擕�iH����*aT��r��1�'S.�E_�AP��{��I�L��lrJ���t~.V.����Gھt�l���2����J�`M���]�o
�p?��ƴ��i�Ң��S[I�&���e�W����nbR^&���:?��Y���� �E'��
�h_�j,�%J�?��p�߹v2�'G��8��6a��L|d�:97�ʕ,9"���G���C@�=��X�eV,��������Km1���$9O�
���D� e��}A�E�i�S�5�d���8��0���=��h�/�\V���]��9���M��ai1�I�� H����|) *�,�l�NDs��m4� ��p�,�"EW����R\c��t��^J1[se�p��Θ�vw4�;���aUE�{�ǵ����d�YT�@$������Lh�����6��,�y���]#�p}����~�wN�X��}�hc��kX���\�,�{9��Y���6�6PSo����!�'��X�o�pyN� �&&3������� d_��D�W�̆�8a�����6���ג+��3瀢_����g��������9Y� C���1-�KM�Sq;�������y�� �u'pmcp@\c'�_V����kB��u�Q� ��,S�s�(�==�B����`b9Z������n�b����Fr�뒕̰�Ԃ�w�	ɉx�0n��A��t���LW�1�)mu(/�����*.J�JD�0i�D@�@�q^h��vP����@R�!+=�]��\,��98�Q�r�9�_����Y�� �bY� � �h'�:�g�����I��
��?	��̦vP[�p�0�zk�u~�2`��5��p(�#'j�2����L��q|��	�>������JP_G�tV��'����R%J�����ebHz�.�:�]Nm��� �8��9���|L�p�󺤏[ʋ���GE(�)μ��A��������A8v��J@�-$�Zr�TQ��gZ� ��A �q,G��gKI!�	��s�Q 7���� ��Ջt �G//X��0�,�B��4lݩ�p� ��Ʉ3�A,��%��,9�\S/�R-��5���&�ۡ�K``�b�Ҹ��3���)ѡ����Ki�%�X��x��(\3��_9��&������dh�F^���bbC�_@��}j��%�� Lfp(��	�M�7��P�� ���QĄ�[n���(\��한���&�;8����;��6�yQ�i-��%'��yq� 
���"��Tn��bH�u�%��I����T�O*�4���}��ñSωd�Ļ�(���P�-"��Jbq*/��,P��o7��|���^)'1є�b݁�V�x/&4���bu<��I%�2ˢZ�Qv6�LpӋ�y��닉���]��!ѹ@����82��^j�T:`%0Pr� (�C��
 ���P��s��'��9[VS(n/�����{�o[~�!r��(�9v�-	�Q�+��-P0M����M�M��3��SV�P�Lć�0l=��0ϊ҂� b ��s(�8 p����HU�R��+��0��ːl�"���.�n(�M����A��%B���`К�.������,��5��u�h=G��� �`�m>���e����噥rjo��,_�p&�ga+X����mSW����V�D�\Bm���,�������&
�E�:��l�/S����$ ����a�����>��4N���L/�~'� UjZ� (��'���YSy�8`֝M�,�#�[�!�I���(czvv��t�J����m:ؽ�fo^ 6T5D[�A�Jdfý��;j ���x�{�̩��Hk�D:#�ޱ	��daJ�R�)ȉhj��<���X�����:{o7��*"�q���$_ ��L��c�s'5R��D�RP���rʲXT�)��#��,lS�}���'t)^�kY��pF��g��r ��� H�s*����	��7@��À2��
���� �A Z�������;���R�M]݅�%F e�\k[�1S��tx䟫��|h#�2�$
3�{Rr<���Y,76���'5��N��H�x�ǘS���e�j?9���'������D������Y!� Q�ΤV�V�9��K�2P�,�\��b*����W<== 1��wo��{wXg�[L���C::~B�=d�A� [yGr~~���/����N���n�i�N�9��S�e ����l�ԩ�d�5���a����0�`���0 @a���<���c��b����a��{6�r�������e�g3֫�JV[q��S��]����2١�aSp	�\�Y�׫T�;���[i6���`�J2��~�z�� &([
?����	�CA|��q����6O�zs
,U�]�Ѐ�g>�m��O��E�[��a}H�'$��٥>lQ���K|8��1t \&9GPr5v����
U��� 
L��ɀ3ak�|
�rb�������CZEQ����L)�~`�Z��� ��@��F�a\9qop�{��^� =1�rz*�&�J��@۷�P�C7���]�[11�bq�e���)K���Y��]Ng�9���Ҥ��#�m	�.��{n��8·��&�p4�m<���	Vh�R�j���m�&�f���+8����@���=�J3��, �B��,��q8&� r|S�Nĉ�������� ��>�z_ߥ���s���.�{���0�wwvEtc`z	u( ��Z}A�ƍ.$\� �l���.�Ͻo/��ZO�(M/,�Ӿ��%�U�&���ɐz5PD�kS�� �x���3��i�YI}�q1,?��N��-g��"�dե�&q�ܘ�I�ɤ�;#�z��:��絷��7�<�����%s��179{t״���2��1�:�F.��1��y���\)��C�@���������2����/�6P�P=Ax2����@��������xRz�XjRj��A&�E�XS��1B�~�(ތn-�����TL|M�	8����D(s�c���Z����}��8��WêЃ���0�Rz6G���4��R-������ ��!-�����^���_J*�(GRi��T䉓�[���b�W}Z
(*	�X����%��7N��l@i,��:-��*�����qZ�F+"��s�q�����赓�p��U6�����$�J,�qPVH��Klpb'垜���s����.�,Ӌ+�)vٛ�\�#��b���u ���[��Ť\���t�Z�ǡ8;��ޣ[��/ѡPCGcܞ���ʡ�~��ؗ��C����_����㇗�/�)i��E�[�� i�-�"��[�k��҉��^X�+[}\K��=~���R�P>!����z0��_��Y� ��./�n���A��,��r�SU[>gW{N�$�bP�w�t���  �t||@悦���̱�>�?��r.m�=�V����;�(���V�>[��%�5j&���$r-`Y���~&S���
��ϴ��M� 1�h@����%&�tu�����V/�R���� �|��q(� ���)��	��E�����O$��&j�Xre��"���ӑr��಍~تj+��G,f!�j���w8�
΅�{{��KЂ�j����vĳl�P�lZ�Jo�bu�_����	b
V����9�T9��k{�M �&����ҷ݇�|^�r5���M'U�S�ݫ�S�o�O�'Z�)7�� ����2s�5+W�`M��P �fY���p��'¤*��z��H��F�k(H+�U^=d3U�8dr�L,8E��>�Aw�i"p'�k(f����؝*ul�ќ��$�����&�*3/����h4��U��C��&�,����M)y5E�AUZ4�:�k�wif�+De��fV.���\޴�XfyQR7󤤱<�W)�b�)�S� �o�>	GA���fa�xb�Q��Z���5���9�^�bhvCv�h0/���j�V.�r�|~��鋢�<�6p��X|�:�xL����� +����h�oʹH2h�N�#�x������z���Ѣ ��E�&�D�b!B�4�7-�\� �>�E(�Qe.@#����a}vi�6��>	�q��"��	n� bn�=ߩ�r��Hb��u���):�:���mbms(-݃k�I�HHh-�X��i�*AF�O�Ԗ5�T	�X�V�.rJ��f�@	
��tc��TxN5ِ���9kLX+d��pB���hN��C� �H@���D[���r��^D/�e0�84�԰~��4��vP"�o@Q
��a�徯+tƢK\]�L�ϿAY\j�6l��"�WЄ����(�����o�3��m:;c?�� "T�~6��}ټ짥<җrC��\���������;�9�hc�](��E���Ѕ�p*�.�s���@,b�,Yȼ�J�
��zq_�k���&}�q)p.�oH�������E�E�L�ԕf�r�Bag�n߾����gN������~v.��\\�9�L��{�sW�g����[��֜�Fk{;�i��=ETk�(���G�T)�w�S���{Z�'I�
I�(���_��f��c������~�18���\�DJb'�U�p��dEm������i�Ծ�B�˓����N�o���?Q��$�6K�����������:::�d��`��p}�C�?���e�u�g�����񛚍k%i3�Z����ݶ��Xu9��}n5�t��xI3����操W_y�k��%�6P�(��
~Y.Ѻ61P���$q8V6@�,-[��˯�V�TVd=Ȅ{�r/Ϣ�k�b���0G#�л,8�H��s���	��&����C:<<dЁI�Ώ����yY� �c}�� ���c-�g�r�wkh9PL�|�6�R7m�D��2'-�I�hM`;�z�R�fA���i0]�Ǔ�h�|�+�#���Tx���vn�>d��˓&�u�Z� p 8=���"Y����V�K�9��9c�,�2]��?�{l�jn$9���5\�u"��
����]D�(W+BK	�s�Ϊ.�KqPK�j�&�np�/�ɒ'-"�/�����k��	� ��(m�c͙��.{ɾ4H�k/�j @Yhq0�?9;;�m:�`|:B��q'�W�M�T��xr��;rD+�H;q�s�sl3��,���7ee��X�YR]J����fyƄeO}_�Im���5��Z�a�ÖYW-e$��k�HT׃"�8�u���� ���2�3��Smm�J�x����s���X����r���Z��O���T������r(����Lm�l�J�\����y�9��0�;J$��9؎�%ͣR�Z�WZU�&�It��c�%^.��c���m�K)QT$d�W7ܥ[��2���|���g��|�8��v��J�J.8��fG�A�ΐs�H�A�y9(U�vm�	�x��q�&�S�Ie\���<�)� :�t�Q���³�2�W_H,j�m�θ.�Z~�KYj�v��h�u�����w&��ɼAs�	���?�XD)��=�����HI 9d@���Ki��C�Y��2К��n���3�B{(uI"���S�L�����4s3�E��o���T�}��X��m�X�:9��TM���>ϭ��KB^��X��Az%��[�{�w��R3���+"	�ĲSU�nꗑ[�Lњ��)c䐚:���6�;{t��=�w�z��}�}�6sVR�CRJΦ4_��L�+9;?������ׂu@ae�%#�._��3S�w�:��_(�%��7������y(h�C��P^2�D��C�)Y�]�hV�/jF��p��Ӛ���V�vK�܅��(]I E���� Niw�  ɫ��+w^	 �O� ŲW%��ۀE�bZ���cz����30��,5����踪?5�;�?G��  q�7�����kPRZ�X�8]2>R.�>G��sS�w�͇�2��J�\�}��ZbŬ٧�׋y.xV����)(���=�Z�@� �x�JE �A1�h\%NG$��r�j����<�o��ɫ�3��`���x)���W��n�NO��j�9��(��hh�����/��f��C1�Ա�n���ҕ�I�[jf�
$L�z
Z/��[@y�)�´ܲYV�S��H�+K;[���q��\��2��u��
�1��U���)$/I6t�`E�vq��h8@r��@98�E�F-x 8�������8w a-��:<ЩR��b�%S7G� �.�e�:�{{1I���/��u��l)r�dR��̾�w2r�'��G%[z0���ב��T�x|s!lYvx ��~N��b$}�u�-;����>�����S�ΈŜ��[̕�0�rq���X�k�%&���}��!B�"~.%s*���:B��`���V��֬�M݇� a)"۱V&Ʈ�z��o��^��vf�:�j<��Q�nA[+�;Oȃ����H=��t~ �S�#t旂:�Q���x�4�+!jr&�?��"
����� �x�K���6o(�.��v$ ��I ����\��8xľ��W���k��D�}Y��E ŋ�^��eZ�V�w.i��u�崽�a����>e�F+����M��o��/��n���Fꍊ�$�!�YǞ�K^�A ���q�"�!��Q�#ߝ�*���|K2�\�H�H㼖�@Ǒ�Xxܹs�7���qE�%b̙s/�!�'gg=z�=w8���s)Zf�y1��e4S�DÓ���K&�rfyF�s@�3��b�fJ��b�����6m�j�Z�ֱї��T���kl�N�8gl���M�u��4�u��1��b	Ӧ�Z@�t�n��q@���e�Pd�8�U�6�V' ���~X�Y�y嗄9b҇��L"$I�B:)u1g�n�b=	D��p$�6L[:9>dѬ�^�}���8���,�:�0?@r��W���l���W[w��}O��YTnb�P���!Bp5u+u�Se����x\��ӶԤ��+��2.Vb�j�Vʚ�`I�r���X�+�e��4{>�Qp�C��B�GC:M��1���s��j�Pe����3vU<��ڏF;Q\�w��˟�X0�Z~�Q8��wt�t�<�ޱ� ��
"������%����$
�d��9�����e��]pB���'��9bQg�`,�S�K6Ͳ�������ڕ���:�WĚ�r9�/�.�Cb%rɗ�OkΝ�Mi���I,O�ɤ��S)@��u�Vg�P[�9����%�֠^�^J�0x��� n���z||����:�� �|��>��W�3���!����k���^{�����g_ a�;99�cശ�ӥDB/��T�� Z.$���;w���[����ޛ-9�dY�W.��ᑑ�UY��5#ҟ�/�K�����E]�2U%�#��᛹-� ���E if4w����F;T��{���o�gr���D���#���*5j��"�M����D��> zh�;��m�FQ��`�|o�	&V1����0�g�|`S)�P�C��ӣh���Q��j%�0�vt��E�n���^08��ڎճ�s.]Q�V՘�����j�����O��O�L�`x�B�Y.+�d�B�p�l�!����-_;�q��Bt�����,�Tr͒��W7K�)�aC��:3��6w�����Ο����sP��ŋ\�M�.�i�xk��+�H�%%�T˿�zZ�����J=�9ŅJ�#ת���r����=�!���ê��I����:�s���}(3*�jă��fƠNy\�����<�A��d���[�` .�
A΁AϩZ�����	�
e0�b]N(W߮Z)�w2�]�?�m̥2`g2�]s�{�:F ��X�2��o����q�~�M��n2�������z3�:��I(�>�%�RJ��p�{�D��3�����H�>� ��D �	�b��N��eձ�:�*}PW�����DPe,�:���	�W����t �d8�}�ɥ�|��Fc �7�i��H�uW&_a�Y����Us�J���I��%��Q�C���y��G�@ ��`<�Ϸ�P�A_�qO.ɽ�j[�7��#`t�]D�ĎQ��Xtcu��K��������^��O��e�c�Nޱi�(��Dĕ�2��N���� �[u�h��� 9>>aPa�Ѫb"w:5��A9���4��}���=�T����r����#�F8�l��VsZ�R	�5I�w�*�������C�����P61C*�=�Rr.�D� M���u������~��/Q�VA%�g@�H5#���l9G6��"�I��fvFǃ�j[n���
i����dAz��e..�,m
���:�����.8&ǳZ���r΄+G7E�K���	�Pb�H>�T`Og�i�]@c�Dir�������2KO�n�ʃ��I��Y ��R�E���������Z��_(I��o�f-��[���a];�og׬n@�8:k@����1�� e �M[���h, ���U=���������y����5]�\1�"��+�N�}Ҋv1b9�M�����ڂ��C��p������}���s�QRkr�qL�2H��ňYqp�������q��LT�A�EGgg'L�"�<@��ǫ)]]_ӷV��DNS*���2h ��H�^�' PfQ���JF�欬%K'��Ź�W���Pvi��+��2:��$�J#Ab)���W��^ڡ�`3�1�9�ʑY�9I�5�$�� 2c�"zwҪ* �0���qć����w�p����m���ng̕�fh�&�<@��ذ�@�� T
�
��� Rsn�ZŮܥn�M�7b:��f���4;�^g��}/�ҿk���$qߵ�$e)����c�O0%��;�)�|pbʡ����d܈����Tx�����^�+���� ���O"�A��w�F8�]�Jsu�dpx��~',��-R�4��[,J�	Zx�r�C�Ia��GՇ�:��`r�6ȇlh��������[�ڷ1_X��d���<֘w�^ ��۝zU �	L=$�����D��*-Wid�֖�|�iCGö��cX�䯜LS*H�����$��H�q9bV��D��3P�@ S�P:ߣ�$WmR�����>�d�$k�5��琄�3ב�R��w@J�J
'��{�����P�7'E�I���d��x��_���25��Ր&�\\�����Z�|pf#r�M�f1lÄ/IEB �d\�4B�1
>e	wno��=[xf�#
�b�������� ُj�
7o���Ŧ�]��R�&@�v�C�bn�yA����Ht�Ya�"=3sHr.�f�i2�)s�[2���5���u�����I��T�z�ã��\��< K�^`JFpT,�k���u��@r��BH�)k[�_�.�#�>J�J(.�Ǜ��|U&:T�������@(YrG5S�}r�x|�;Q8W��O��,}O��!�C��z�ۡ
��;�����r �(�;yX�ut���I
GI`��q��K��dp���ȱ�J���]@���rE�GS::F�eHSS�-�ߥ�snI�a
�kym���r�	m7���:���2�'��%��_��A�ߗf@
�}#.���x��q�[�`h��i{�C9�v�m�A|�΅���0ӹl��hw3NBH@�4pl��M�7#��V�+�
���R��E�s�_iD2��q-�S �!�t���Vu���:J�e���`�:���
>�%|r�T�N����&Pq�����������{t��0���y���;s����ʘ�2���(%rS��{ �M
6�g+���c׋�w�7�������!Jh��ug:��"ZƗ�6�&ʟ8�4�QjbSS ��v�H�Eړ}:K
RA�)D2)U���5K �;�����_Eͦo|mjI��f�����O�b��v��;=ވ��*}jD[��$�ν�(�f^%�쥄-,X�K�����6-Z�I���r��A�Y�
�,!b~�}G�8'/�W�`J���mUŲL�Q��\J��{�{F��
X�7 �ŕ*�m
�f#�ن�i��8��x�Y��A
�*5m��$_l��`�©* f@p!��`*X5Pix&lu�k̹�����>��TϘ��Nd�,Bb��5�3��ҵ&�g*��=_��"�����S,����ua��
��$]��kھ�E�uM�>;�K��)!����*�2�mp������%��~�5��y��j¶�G �"��T22酷O2��Jl)A 
�h@)� &���(�������T_� �Aʦ&҆�Fh�6�u���� %Z�=��m3SW�ծH��M�2�ǒ��M��:��J�h@ڀO�y�J�N�ǆYZ�����#��lU�v���[:>:��v�4�ˊ=t߽}۪H%]]}���k�N-�|��� �nW�z��N����ﲭ����X�c-�*��#M�Yd�| {����β���C�3�'�2ԯ�vM�y� %uc�!(��'�}7���l�s@ARNVD %	���]U��й'���ɘ�<�|�������:99��n�we�h��F�RӒ��]۶{m�,�*��c�8����)��Ҥ"�l}!�;$J䋝N�cp��v��A�X.cN}Pط�IUA�>���b0�����D)HD���8��T�X�p�C�GK����2x��Y�G�k�5��	=;�h�*��^�_��N�tvvʄ.)���p���@�"M��={����)�f�n	9U��[����m��̰};��=���9��SW��S6�t\�����{0M���t��ecci�@)J�M 	`�Fu@�J�{���ZU#S{�p$��8�%"2�T���
(>v�1g�?�Y=�p�U+�����1|�`�ܶ�/�NZU���*� e�� \�9�/��ܹG��ӧp8'�CNHA��-��~s�����Ior���@��{��Fm����<F�q�^�P�T��q9�xz�:�dB��`�B�&q���{��!�
�T½�'��f�HB�q��I�**?�z��K�b�fB���7�؏آ#���$��L�Yu G@��0B����/��ݻw���~�2!��k��� �&5�>{t���
�A2�J(=gJ�~	%��dF�ڟ�9��	,s:��|�L���2iGW��ډ����2w�TR��Y�gx��7E��?Ud�H�قC�����{>_�D2�-��xJG�N�-K�x.�^���8?�b��^�����0P
h�i�����H�h�D%,I� 纁'��G5vL�#K ���C-��J�����쫵�|I�Z�9i$�?u`c�l�;r����!upD:��Z��WR��7l�P�O���趏Ou>#�N��#'H%e!ŞPYpsc ]A�0!�&ttr�eI/ @ȳr|B�޾����E�u�,�5�&��)V!��L��ʮ�����Rt�q�T�&\�ow���Jߵ7��1S���v@k����)4�e ��(� �����[\hz t���+�P8O��� ��˝ 0�V.qEA�W|8� [xJ��Dg4��$�� Y{Bg�	��b
ɲq�������/�0	��T�HB�9??c��e(�.*�R2�!;���W��o�C�/��gV��k�@���l�1�v���E���a�g(�ۆʁ>d�����QIZh�Z�7�[V0xef�3������(��?�T� *�ZP��Vi�|�t�jV�4Ѯ� ���F���BKj�=K"�鏿���8(�!��՛��Z(���@F� 'Ҋ��\)��e�kb��M~ ��'y��Dn�{�u�g�m|P�t���L֗�z?��^r�>��}�!>Ʃ�ȝ��\���'�< !���'�L�N��NݔFu[g)i�b�a��^�Rjc��>���������?�����4�3�u ��,�H�}C��k�R���������\��d��bH(2 ��Am����o�k�*�йA�I���&�e�F�6N�1����{�g(f6Ns��7*T��*��H
]�C�Li��J1(���
\��X�d�:s������z{�H�y��)	9��]����S��LPH��M��ӟ����������0�9�$g�R	֟�s� 	�0g�� ��b�������/eO}<������a�߰4c���$��`zh.�⤩ Ѻ �*�sݝ���g(�9WA��N`� (���R��i:���F(�f�+8�0ĹD�.���ǁhJ&rTsAJ�6dAc ��obu���7���;�P`�����h��rW�LL������x��~������O� [�$�Ƶ7͐��ǵ0�C�����	�!ߗ�߉Q���/˿H(O���O�-EpZb@�P�b`�̄΁pȵR����U^t}�	��,�"�Cժ�8�#Ad�0�,�L�G�?��GvNC��/_��o�}>��L �g���^޲���v����I��������Nꊂ��As�X�7Y|�_��>�I�K>h:�H(='���U�"�<jX��t������}P��� -�`u7��i�5�t��g!4�(a�V�s)�1R.P�jR;91�h��t�Q��q�׭T��cC��|���ӫW�2��b���>a�\I��o�������W���c+��0I��JÓ����l�O����Ѷ�3�Z���y�z�t��ԏ�B�	����@3��{#�i,�H+�2=�C;0#)�^�f�O5	Sx��9?t��� /,@�/�����8X�y|i&a�9���H��cX=��(F�3&dQ����ڋ�-�Ƴ���=A�ʏ�N���G^��ۓ��4;�~�+�B/��u �D_!��&2Zp�/���ځ:�M_�\���x���R?���Wt{sK_//�XpP"���'��̎f�rFc�Q 9��LJFVlIBM |_� ��E\]_JZ]_�ti��Zd&�o�s�T|L!��=������`�}���4��e��r��N?SS�Ο�S>�8�Vv��Hܳo�,�Iͱ_��U=I]kI3��%���ԛv�F�J�t�����u-��Xy�{[�Щ��@��Kc7V}�tl�.0��QV�DH&Ӻ�N����� �u�{�����(����U�ޠB����^�Yz����F�K"(�?���=_ eق�޲�c�n(�! K�&"r��"H'����y�S��4ϼ�~�5�(_�F���_$��2����Y������Jw]��y��}Cj0��cZ�GT��a�a@�8)�����-�$����b�6֪n�.QM4up48�v��bn�����<����0��K�^ 5�/����T��N�������v���e4���.sQ �,Ϫ��������$G����N����d� e1,��Yq.X���<K ��<��yA��d���D2�����&��
����uD�U.b��� ňO��h��d�p��w�&&)��Ԣc�ĩ�ҵ�0��Q'�L�3Иlg|����p��w�����62Z��`%���(���,��h*�)� 7�qt0����g+��~���%̪��4g�^�_���!1�����H�_�]��s�@I�ڷjQ2 "�FyE2��L$���@*�z�[)T�+���ݦ�;��L� ��:�m��%�ݲ���FuS"dG�a�	ڳ�]��&��:'��g-�,yY-�#��؀W�O�U��o�@�sf�����Wl�"�V�EcM�S	��x�՜=aWՂ�/8��W�sr��ի��&5�D�YK�d�@��[ϱ���M�������g>!�\�S���|N2	"����~�w�����#�u��Jx}χ^ ��7V\
��S	E:d�yY�R�$&���m�,k:::cB)�t�x��B����{��XAz�%g��#���ŝ���j�]����+�����6��W,���X0g2k�����%~'���0��=:�q�Ig��+�|G'M3��@	*��/�;���U����v<G�(�\v�a��EBy-��� ���4Se��V�Y*�Ѽc@99n��i%�e�Ǻ�/u���qqѪ-�<�N0����I �ѿ���@>����ԃC�|q�L��0T ��$5�>0II-Y	�aI���݀�Y��C�?��� ���?SI�y��熳��s�w�ǵ���Cc��	��\O/�'m�{�t�'�~^\�F�˗�N����)���MM����T�8#�Oi������L�ZF�dޯ�J�j��?���}��w�>���?�W���e��\r��ϟ?1G2o���t�~R Q�z�O���Ɨ��%b�	��*}���{L�������K¢�jM��^����� %}��\2�Rsb$ߤ�q��Kĺ
q�O�^�� > $�IHd$��Փ�[��  �l�y��s"vN$���矨(�:���?~��&��@��:��@Ev_fn�:�"}q�G/��2��g��&��:�}�M�v�P��}�%�kq�J(�g�JE��zy�(�v%��Eh�c�e	��o5;(�zv�bd�Ë*��6�Mq��妳}T�hH 0�6�&h�¥*Z5�c��ڇ�q����s�|���77W,�|�����4�����5Ma<b߳�iT�I�u����wVg�~�>�v
�?z�O�)�S@�p{ %U���BO���/YL՞�
LО�iG����l}?ʭP�L5Kx��<��Ņ�&_�~�Lj��A�
���+z�.�R~��7V; (Uu��\]_1�������R�U@�:����;KޢZ��6�.�ɒ��c�F�d�!^ ���Kj������S��7o駓�	ި�X��]Hbr�|�*î� ٰ��k �f�Q��l�h���`_��CK9?� ���f����Lg� �8�q��~vSkD�I%�˥�>���dL�,9���������߇H�5��Hn����SW�����b�� �8a%�wH�Cn�)es����ds�G�l%��R��B �+6%0P���-�|j��2s�/�3NY0jF�ItӂHXx�B=�4�mW�UÃa<.9?K��S_���w:���^E���P� ҧ���\�=�8����B�7��B�Vӷ�:ҕn�a�mb�9��� Ŝ�,8�V+A���Y����xJE9�ׯ.؁�4V��Q7���,���+����m�= ��O�5­�������/�1�: &Hba*��:���G�95���Y�v��vƲ��!I�ߑl�'�oF�M������T���:�a�"� >�\���G�:���]�u�q�^��O��������'�h�ׯ%	9$��s��� W,�u�J, Ya6F�$ ���D\H)�?���
���G&c?�Ĥ�8� ����,P�V���2�Yl��w�K�D|��X&���;�.�j�,�K�]�eMBY?���rdn����黮Cl�PXδ���.ė�Z�Z$�SuE���
����ג�~%���I�7���8�.��`"��j�I�nnoB�/���_Tl��g�M��|��@�c�:$޹�c�5�ha�9%m� �����i���.����n	���9��e`���CH(C�������Qާ2n%��L2��BT1��� �r`�	��rI��Q�^�eB�7%�N�r�֖��D\��k�}���ɉ�`_�K���|)����U�C�lɎ >�U�`���ɐ�>WW�\�~*�JF�.X�޼yC��*����o�����_QY7ɠH�8�fR�|�ΎO�7�?�v��d�7ls_	��;n���������n�x���D�1@A*�G�0� L�i��;�v���Y��6 k�0�3�&OJ:P��֌KG#6oU�W�ްSHT����^pG�IV#�ng�ԝ�����H+�8`>-���������]������t�/U��u؊�#�Cz�̑��C��tT�M�_�������L~O���?t��J-<�5%=�HT���H$���砐J��!�8�Q��f�ݒ)u���e�n���'����aQ
׮,���M�>�p�� m4�R�5�	Z�1PX��H��Xv7��g���[ONO�V��ot���0�{�������*�+f�n@� (�\TLT�ӓS�:�P�&S���`D��_�Z6tv����{K�������_��کG풯ջ����A
�
�!V��4ib"Ib��H9ݖJ/��d;ej���z�68�q����$�~��Bgt������t'$�d�"<�2)�yW�!x�:񼕠MI{!����m�N2�5⒵*�q��J
eŁ��Do�v=�d�i��)u~���輀I�%��So�
(I��-��F&����&���|�����N)�r~��K\��H��9dć4�@����7�:�	���(���V��''G�~��}���؜�
�z\�\���������|�lϵ��A���s8a'�: �nąY���t�WB7<��G���O���5��@Q�Dglu8ty�
��8�ao%(�r1ަ�b������!�eMC3+�����6շά?�7"��+����.��J�^M�ڄ��'�� (%�TDhjϡ�`ߏ�]8Ua9aph$zעvE��
 ����.I��$s��H�ܮ+�����4%#T+�usS�z���U�X���X�p���2�D��h���nL_\�����'L�"b����i�}��-y1чdL uq��Ѣ�$*5�@��H1k�m;���S��=����Q�eHd��IMl�ScR��I
��Ʌ��z]g�;L���g�g!�EZ@�#/�
�#�C=�4�h��a˕�Д����:HU	����l"}�vBK�$�����#�{Ʌ�!�����3E�G��:R=~�k����_�����,8k�$hbއ5���`�~�yS</l�r�4���M�NmP�u�����1���[ߏ��#x��EUf��	4K^���R�u�/��w:��y�@�c�=;@A�9�*l}��;��gĺ���D�Agh d
��@��>��
0�����3vx������l5	�n����\�G�dKaw�>�	�G� z�u������ӟ��}]��q;s���߸OU/��
9.�! *�oC|[��Ε����� ��>�8�|�3�;�Q�F�ȼ�;��^�#X��G{v���Y)¬Qז�b@W2i���s�¹`�|6��3ԗ�kb�-Q@���ēt�R�D(;���I��w���(;�@AHGXF�2�$Hr>
�7 �Oz��1D������Jŝ׀{�2fCb&�:��O�r �
��Ʌ�O��X���t�s�\���2@��X|#�3��=_���o*:�X��f��+�&l>T�c�h����l��R�����dg���eɄ($8���S?��Z�3��f3l11/9���/�/���Ɠ(�2ؠ#â� Ȫ��|P�K�(�jjZ�X"�n8j��N�*�8ޔ,��<�ޞU���-D�ڽ�}���p ����+���w_�N�c��>�[����z���[���̝~m�-7?
�����&�R0H4U��
��a��	�Α�c���k笂e�T8�v��1��s&H,͵o8۽ӨԊ�s%��f�(\����#&EX�������_Y�@��W���z�횫�z \pj�� � ��W�}z;�-5����A�lA6K}|ߔg��<�pH:y$IŹ����c�8���I$Ū�|�����?�f�Z�-��k,��pqGޑ�#�������:�T����+�
)<^�x܄:���7���d�/K#U�H]]�
��%�F�`=K��� m�09��@��榕`�|�&��:��(�q�F\�����/���4H;�y��2�s����ЌN�U]�OK������)=c���$�2Q������!1������~�?���yPRʳK<��o�W=b5yK���7l
�R��@�b0�W@J�Ι��ҟ���l������I�G#>�x�.���b߆%�{�L�NYŁ�O[��x�]U5R�CU1��QMp<~�"t��V��zA����z�"�+v|C��&xor����J��0g�n���)�V�3)U
���yO���>���q�� ~���_���ڡ���bT�;���`s��\�b]����q>N�LZ�b�䨀��U7ZA�7Y�1>�RZDP�ņ��	�t��=�X����֫o�h�j��	M'�Z�4�-�����|V���c��z?y��͏�u<cN���P��n�m��"�I'��d�O�,�|lRU/r�9��Pe�Y�-�L��E��+����-b�aG��k&Q%j�"�y�0CI�G>���Re`"̅w9q���԰�˒�S	+�S�R���+:=9cN���~�������\i�+�/f*وW��m��T3G�V������&wܑ��n�@����
%��9YM��QK��;��p����_��ڡ��7���K�~�\�[���*�12���oWJr�آ�,�!4�r�Nd������X�@L�ҷj�zͮP�l��3,N _��]_#����Yd����������;
�s����}f��Ҭ��.`lO��Y[�>��x�1AѾ����h�u�T���@�E&�������t�˵��c�C��ffc&M��`p׵��T���ԋP$��A��U����1�N�
 5��¼f�ƫi��,�$�ٍ��v�8&ም���lA>(�I��,�lu::�һ���G��9A�^]���&Wڎ��mЊ���﩯�>[P $�>�پ\��ۥ���+�i6�sq�?�	ll�0����`�g��Ŝ����7R�4�!X-�<�y"�����:�&5�k2VG�Z��0�Y���cqQ�v��loA�>�s�2"���������s��].o���ʝ_�fIW���W8Q^�AM�Q>{w�$M�Ե���Y�z7;�@�j�:�1HX�T}6	��!��	������[�B����0�p�p  ��&F�o�K2��}��Jс�,&	Y�F�jNB!�J`��*����Dbi�i;,F�������j�ӓ㠊-W�b!j�AuC~��Y��[�g�좉qC��L�Z���5�7iT��g+fx,�#�׺�ھ%&:���PL2��ũO$ �U�0!���'�֐l�a	'1��\�ּ�^d��M�� O�l<��6�SWu(e)ޮ�����T.�/��չz�b������X���6�D��L8���LME[�A���	�z��DrP"�#�g (����f�(%�ķfYj����j}�#+��̙Ksv��:�r���x(���ME�ZwX��GU��dvf�Y�o/��H����Q�^]s)���ؕ ���M����)f���3oC�'u;�����*�Eάl�#����	g���q���=�pr_>Q�֮�bԲ���Z��L���u�|V 4Ɨu��}�2�41�>XU���/~(?�u@�cVd �`��¾%��/҂�7Q��N\�^7U��dML���Kʈ�k@�P$����x�֔bޮ0����zo�٪��Z����А,��^O��(H����M ��e�x-~���c-s���ջ��#v��T"��@ɩN#@IA<%fӔ�q����e��M
P�Y���m1>bF�ĬW@1n���;�)}�b1Einwuh���u��1�����$��J�;�iȥ��NM;w u���l�.'�ٮ��p1g��˺����<>�%�ߓP��{:�����㤅�s�4�_����ܛ���W&�+��1��k�F����f�:gjF���ݮۖ�oߝЁ���N�>��M�hX"B �Js��R��M���4m��16�|t��s��#P������;���ۡ������T�I�,p�d�iԯ��K6�p�S�W8�v���N6F�"�=�53��9��������N&�<����_�cۡ�u�̆��{�-֞������1���6�������+�D�&~ǧI)�?L��_�f����vI�~߲�����# �Aq�
(3�d�0P{�J���R������ �[-��3�����o)ײm� %s��k:�7��J�nM���9sҔ�$��qlԨTҽ	&b���1��(���ٱ��u0���l�#Z�{��$t��k�b��d��|�{_������_�9H:㭩�<�m6���p�m��j���e�v�z@*�P8�L��������I1}�]���v��8���)�`�#�H&�`�&#�;�M�®*Ϧ�'Q<dd?-	�>*�>Ι�?!�a���'��ɍd�R���f�<���q��x�¡|��ז�iO %�>0e�<g�$��;��L�������N��cɺb��x����1���W��G�J	E
,&-RB|�&�rP��s����Y
Os�@)�@/�c�|�;�z	�f�-� 
�v�>�̠�5��K�ڦ�tՌ���ZI��}���n�}���C[π��ׂtBq ��EA.u�CK�k�A|P�Nԋ��[:�u��
3���0���]������"Z��w��=����J'����{ Ż�a��L������ QU���.�J�D:x}>2��cG���Ռ~���1�.�s?�}��/�/^ �)4����YM׭�CS����C��ݖ�6��<�a�Mw��n���-���p>�Ԟ-�0ωۄI�>�6�Õw5o�T�pۦ��F����h�M��!�����H(���,d�[��}H��I���=;@�bk.>��@���BV��}�l���Y3�����GO�UG�I���j�6C*OpG��~��{}��*�������E�OE�����Z��
A_���M�fc��{s;���h��֗^��m�\��zH����/V�����(�hm_4���"}�;�q(�c��F�ޕ��w���_����h��ssQB�r�E��{||�elc7\S#W��ɝxZO@�u����C��-����ә)L�Q��N�l?B��f�dr0��v�t=n�����j̉�|}*mB�'�H(e+�� Q����c��d�>r7U���)�L�4������ow�?(]��
Z�I���>5�X����	�4�tT�rlٕ_���'�����I$;9�|��_A��ۆ�1}bpV��s~�Kֶ`��x�T���I+f	*�F5���v��3���J�.Lp-`�H(?�E)�g�(��6����*`��t�;=3��O�q�}�-M�9�ڶ��Mg�\E��cl�&��h�KtSg!���:�U�D%�y?B�%gN�ƹ���1��قJ���p*G�?b��>��:��
EH��@��(����|X�@�mRGߌm�E��byH3y��l/��m�r�Yp�߇����a�cw�}Z2�>��~O�sM�Ο[�#%JmKvu]ߎ�O��;Qu�+$�h�$�4hѪ�D�D�;��Q��e�A�����m � 8Vʕ�zLó������"d]U��&S����������3��}����k
(h.���"7����I���{���y���jQ�=ݖ�4{�	�O���y����P�'�����(��E�����#HP�#�@=�U��YNl���ƺ\M�]��0Ix�xN��9-1[�)��� �|�����P�,|P�t��ɲ��d֞l(����]$�]���c�r��u� ];3��oݿ�#���jz����{��g5�Ц*�.ު$����Aݣ�?��w�IRI����'Ԟ!�t�����>��{w���]�_Ϭ��7^w�5ص�䞆���I�|����{�ʏ`]%ꦕ����M�/�{HA~�wH��+�z�zs`k�srٵ�o���.{Fw|�$;S'_\�a�Dڦ��\��,]t�k:�5I�����������ߌ3h�E��K�J
<���3�8������-+j�<�m�P�Q���lB~���gh���`N��a��\��ƚe�O�;�w��v̇7��_��w$練[��%&.EҹV$�=?!�_ ��۲t���]ǫ���M[�����]�$��˘��kc_ۧ#��k�w{4�v�U�H��j���.�v���>�t�۵���6gӧ����K�X~)�XLj��['�
L���c��#�@�[�>��>Pq�7ڦ����Z�m"`� ��fV���Mvf�.�V@y�u+Sy(IRM[D{k� >��(����c$mW\���J%]�o�l���vZ�o1�Z%�>ۛ�����L��2n�'�J%['$��X�Xqq��f2�W��K�z^�-&�N%������,&�I��!�@���(�^�}��m�}(���N�T��&|��>� G�P�&��>�w�=-�����������҆�]rx��"Q�v#�4.J�͍:|��D�*�tT�.�K(Àҵ�p��-	��s����A��u�PФ��[���4�Z�(ϭ���G�Ǿ��'�� �R֚�7i�S�1���(�B-{2w��pR�&�����Ã�����N�^ ��߲l��.�ﬁt�ᾃ �$��IC��F��ξ&} T���4eA�t�_Ϯ�I�ޘ�Z�T��J�暟^׾,="	��K�^ ek��<d �O�Y��o��]�C����[�n�w� y� ���xY�%�JL:��� ج;��R�j����l|P�Pz[2�8�����!?��;%�|���bV޳� (�w@ɬ1~(�y��`�Al��<�����<4(��ӝ[�6%``R@1KO���P��rڿ��j�]ҡ�@lb�\_���l�7���w���j����(�x���G�ۦ�{{�F�D�^�L=@ ��Z^�P�`�Kg3M�Ʌ��!����2h㈜@��%����1���%̿f�s[ ��?�Z��|Z#9{}�12����������>}o�,G�Z��y���(��1ˎ�Kͤl�U�����m��)�{��Z���C���K��'
�r�+Յ���I�3�Sua쒔���lM��K���[&*�obG�i�y��٨�$��,i ���6��օ�a�g��7v/��7J(ݮ��x���횿�$����P�sj�L�i˓+��&��%Ϡ߿$V70'u�}e�"t�ko*�_�r�U���r��"滼\����ɇG�1���4�i�h;����a�U{�$ә���:\��ZY�0H���Z��'�R���"������3�Ǚ�J>&�iJ�t��fΒ''@��R!�.� Jt�$�d@�\�Xr��>[h�������Ǯi^�(�AT�wB��J"*	t��|K0�m_Y��A���A?z�]��S��w�� ��xtP�Ih(1�U���8�QǼ��ܕⱻ�U!���.���6d	����A����΍���f��<sU�������ɀRN]ۀ���	����?�(��+�n����Yv�k�U�(]�i�dEY�_�@
�3s�|�e�b}'���{��n�蹗��'�:3��@.'�:�r���`�ǧ����8�ɠ'�LD�~c@b  �#z\�	���&@R�q 8�I1�7i����@��"�wz��T�!<�]�{b�$���M�X2���s�6F1��(wV�vj^�d��a��	(ڲ�Y�6;t���$�(��V�h���m���H6��M��E�-�)ɹᒼNs;�HJ��r#�e���O�!�@�R�ҽ߻���4�Lb���g�&�x�o�$��X�~mkm��\t�����V�v����3IN��������]�N�� d��DDw�ɝ� ����k�K��5Yti3��)E�:����JF�*]Xb�F�c�o�H��;��k�4f�J�E�C
S��V�gj��v�=�)��a0F+ͶûP6��ᤀ��N��*lAE�u��h���p�Ch�P��,�
�A���|���AL�{�W��_�)lɈ��
^hʢe�E�D�Ґ�9�Ag�*�lS����K��h�"�9\��'�^_����]v�ܕ�>Q��J(]@	�N�ǴO�s���m��	Hn�����R\�S�T�y�ۯWt(��
�)�|�-�	��Xhȋ/���JS+)*M�
��J�Zy�Qک�,m�}K�U"]H�FK6�T�j�'ɬW�����vb��7�K\�Z� �
PZUJ��jn��օ�W��6��P��qR���ͺV.j�36�����$�h$����f�xx���g(h�'�@^�~��YͶMf)���$-c��'�W�VMJ~��Sg�s!��Q��M��Qщ�TB?�Jx$RH$�'�Zb����|�H0��Bb-�b�(-8��l;}!�Y�eF��[4���P��].cݿHί�Ib*�E�JP�c��Z�B6o�)Wk���{ծ[.4�C����&$�PQ��a�e�7�N6sI^TG��B�MOh:�
�_�DB�MTwR2���q�2 ��l�k4:uTNŗa%>%�=ר����G����Rc�NHK8w)ڒ8_�3b�+]r�I�}W�%(�}��e���O��O�>����C��&J�XR@��X7��i���x��Q�<�� �P6Έ��YuG�h�}�f���F-	3�j-;�Hj�����YRCY�YooTZ)ˉv\�|��ŷ[@���J ��"�����8;U�bA�*%i�ZoF|\���d�u�lP�9�>-��tX�ś��}�i� ������v�c�y(�{�6	���g&�M%�v= Ŝ"��R>����B�g��q���P� d��I�[W��r���#����W!��h�e�JI<�?��<��"��T��:8#���h<�Z�����c�w.�-
ٶ.���H�Xv����J�ͯ5v���Q|ƭ:`�N���֭�{k&�=��ׁ���f΂;]n���8�'9�!�g(�10����ĝ9mig
n�e��ͳ��(�v�aR�Z�ݢP� �R�z�_�  �JY� w(��ʭ�y
�	�x��h:� ,5��ǊxL�B���Y��H��"�t��˯���c���}�O�S��C�g("�"�`�9���">dDm�����I\��ꈥLf��H�Y���P�J=N�@��)��@�/^�1��g�g4j%�o�����޼~�.o8��j�
z;�urr�ǹ��iE�����:�p<��v��&�	�{�����}���noo��7'�X+�Ā.�t����:��r�vTOT��w���M�H�Zn���}��f�7�G���\'�gѠ�=~û������Nw�.�t8�����x�|����c P�ڿ�	�"���Щ$��[u�:���E�J���F���Jl�������%]]]�۷��ݻwL.�vY2x �  8�ׯ_�������- 8������f����>�����>�j�P�����,��$��?k��	=�ߣ���D�	Z��A�k��)W����Fl3ޟ�,=ߩCj�
(�:�,��Ѫ���lU�.��c`�M��#؜z���-��(�����.R�(	��̉�hg Ȩ�߱��2�ٯ=�===�N�T�I���W-ȼ@��i6������T�����L�( $#Pq��������_���:1k�uق̛�!K�gO?6��S.��K���Foh�#��f)���d��`9ଟ"����:>��{��6i���W#gS	�Jk
�9�p��n '")�=�R�G6�sx�E�df��������ӟo#�2�-[)���.11e���`?�FX��j�F�G>�?	���p�B-?E)L�l͡��r�T���	��\�鑂�)SH���ի׭��-:�Z����˗���W���5�1d���I@��\?�ak}���TYI��UZ�	���ٻ�Ȉ����D����h��Վ� ���^��I'h(���^��Eėx���H%�Z%���̥�����nj�r��1#����	�}̦eG��U+�v ��6�/ԎE+%@e����aid6��j��U�}�R������9/bq�z�&l�m�Iq,������}{P�b@`��x�>����Apٱr�dm�����Y�@�N�J��A�AZ�;M�n<#���QGh"��Ʉ\f����`I��R�">���ź��3�h"-���91y��%��k�/�Ǔ����Z52�G�Ck(F�Y�E7�/��x�5K ��x�����]�f5��AU���bƪ��Ǹ<n��\�Zu�Iӛ�[� !��`���o�xfW����J��|a�i�x�j���t}sM�I+Q��"�g�k�j�oa��i-p�G
�K^no��o�ɐ����招���-�ݶd��&����P������8"�9X���@�42�9��Gv��0��+�/K�cM���;������X��$S+�Ղ8�b��D��g�e�n�̳LFb��A�k��^��(,�*��v-f�q/*�r}�P|�_ܜ��[� < �Dx;���ɐ�gF�^��V�����+V! *,�E@Z���@1����@�����-HM�s>��ǚ�T�h`�n;�j�Ί�\_ٮ�����Z	R��Ӷ��zV<�0_��m�������	@�X�H4H(�QOq4�P�Q��<��+�;�z� ��2��=���:���%~��*ME�U��E�Q �d�Z�P��:�*�
{(�u��B3���X�,��ci�~Dj�"3�7�m&��Mh#XV������A�x��e,O�X�,�%����,�&�+�uR%� �>R̊�p ��M�D�k@$>;?e��Z� t��*�ȍ)q��d��{]/C%�Y��K�M-^�M�j��U�J�*�����3����0�-�P�"1s��s��U�	Ow����ʷ�[����{���k2����~*F|���>�Iv��
�v����=;@1}�bu��� 
����+��N]�W�J3�7a2Â� 7l�)UuixPO&0#�	�0 ��!q�:E�j.���B�B
��n�:�Pu���ǬU��,�H>�q+�H�'H&1�W��%8�)�7_�H\��ņ�����}��	'�%��D�ci�"�R�r+U8���k�>�.��XU2SmǊh��.��Y�g�sɳ�.�e��$��<��� -�i�Z��=iK�-������J����vN���ܑ��L&��tr��1/�������\3�"ͷ�sD��.����E{�K	:[��m�q"P��|=�qP�77�a[�Nl���D��S����ʃ{�u�{<M���k�ݧ?F��qۼ��(Gǽ��;�'wP��������-=IR�cP��� \0�8D�,�tŠb��Z���o0�~e��իW�~K�V�y��-�	 =@¿c��$|��Ƿo�آþ��1nUx��Y���}�NBL�p4s���x؜��#���f��2���q(؆%��,�[>(��֧L�Ғ���ι�<h�\��;��N���(����ɯdPȝ���>��k�����[��}�<
���`PG@����R�m����I���8�)x�G%z�x,d.T �E+y ڷjUH�
�dż��r���lE]rُBy���֑:]M4�:�iX��%/T��lv���b]������� g�������K�ў5�t� ĩ_
$�E
("%X��Z�}Eɦ\ �HU	x�bn�!5D@Y
���Xp����\n.W&�81W"3�dhk��+8�D����#u��-r288�R/t���?���2�j���������������!e�T�)���H�x;bP��(�U�@�pVǶR������	s/<^Łα���b{j����Hx��
T���a%C��������Q�0B~[o��f�,��A�=a'��\����5y`��8�}�����F#��mQw8W���Q�RՙB� 0Υ`���ݵ5.5}���O���*w��9#�z=�Ig�˃>����d�eJ�R��������uq+>� �d~�:dj�3jJ=W�v��˩S��r�z�k��n��ҙ�c�a�(��?��T��y���ã�I$�%e����_���o��{��������(�U!YP,#W����
��kދ���~%��VA� ���G'8�k%���c,iz���*R�F����8��{�/U��jz_����A�C�k:��J&��>��DЊ�q�	Z���zdnܶ���8��i�t���x/�P�K��p�e�q�h�w��<n�S��:�`���3#AՁ#� ^ŌL\F����&����m��4t}��=li�p$�e�s�?��)��<�P~В���X����t���@@ Hݴ�jϓ�!�wF{6�{�M�[d<��1��v�Fh���_��4n�T"�M}e��f12�����(��	�odPU���d�fj�|�/�@Ŋm�E�8G pVm�H����>�S��	�5��3�C��R�S\6�ZP�(H��Ť���q��$;m���̴�f�OJ&�P��RG�m-5?o�P��U;*Y�g��ڋ��W�^�D�k�k�p���a�y� �dDV�8k[�N�T\�V &�E����5}����+�Ôۘw.�ābې2�"Sqhj��3H��*��"��<-����蝫���냲�m�;i_�	Q�ə7 ��^��.@⨆.7��Au�I���K�=���d�*�o�!I4�t��n�Pd��ݵ�I�.��6�!H����ba��Fˁ�t�p�s��1��a:F����t�{��s�j$��b����c�M,��U�˹�ԑmݱm`�2;>�����$��w���׎a�׏O[�+u�0�{�S�Ԝ�Ã�LJ��_�=;@�f:h(�̳��x��@�U?�r)�:YG7v�CN�jI���BR"�~ �Zp��b�pf8�OH9�(S��`A�<�b�滴�%�N5A���O�E5!o6����c��$2tn(��,��l��^��Lu����Ҭ3�iQ�25ɩ�(hjMwЂN�le�qPGbQ�(Pq`�1�"�Y���V=JT]g�8C��;.�a���~��sV�㻰k��I�	R^4Tuq����{��ͪ�sokRT�\!OGb
bQ�[ߵ-�-���A��QV��:�T]���'i�@{���a��D����	�rH? +��� �c����(�@tu�Mr���]���]
����Z�vI=�wТTv'H]��R`���fD�΃WIX&���W0��~�h%	U�� h8U�&j�c�oD��ߒ�J�K���+�ʒ'��Z�:����ꂉ�:uQ���Vi�Ci�(e�2Q:�<-��+�����5ig�:3�d!��/�z�X8�(HIꂣ���Z�S~�4	<K��Vx�Ƨe�@Y�u5�=ߤ$V�P����C��F#M�Pяh�1t(�GkQ���Y��k�V��������(�����/tq~����nФ�b8�I����
uH;[�b���Rm:+�͕�S	�(v8N2�dy�T7��0��s�8o �9N,����dN���B��(S�
.�N��V�5j<���	��B"�zJ-Uqv�ޥ@�n��m&_3)�����[I������b���gj`��2�i����{f ��a}6M�k5E�+�$�fi ��1i�0���#��! �����Dh9/u�/��:�t)��>���G����쑒R��
�eDo4�����{�)7�O��E������`�9߫�b&��"�`��&Q4H��M�k��k���#ݡ�@�i&���ĳ�� M���(U��,=�J���zٮ�XjIN�d���0�БV�^RW�Kk/T���bP�͂"]��G~i�@����8 ���t����{�Ɉ�)Y��nB*���g�N-4]R8�D)f�G�8:�)�S|V��W�v�L#Ӡ^��?����͗Neꉤ�\,V\��^�~�9T����uː��U�'b{��+ �5z�\ҿ<���J�S6���c�h��#���^�0l��I9�Nk�R�Fb�#ztU �8�l���jc����%-��UX����=��fϢ�{Q �Ck/��ӌ������Jg����:���1?g�G<��g-&E�|`w54��ֈ;wN��&QXgU�5̴��˜�d2������`F�����cԠt �u��]kIGBI�:h�$�{�	�n_Sjn�zS�˹�]-�!�5��'��M��pu=��\�h4~��f��[Tq���Ms��Q(�� C�דVjX.P��a;8��]�[!v����U���$@A$n��,eA̗�e+ⷐ��Y���#�l>���w��T��Ok|$V�Ae}�B�$�m�T�-�GL�λ�K{�����Ј<�����3)A<^��i�H3�-8�+�#T���@!M9`	���Kՙ�Qg4�� ��V�+	(���;n�O�5Ugh�hݑ��k�fMmr��MQ��L��6+b�u�W�Nכ�#P{��f�� R��/B�3�������'t��䔷���s�]��J ��k��5F�ޣ�cQ��HB!��Y����-:. ?<��l���g$��}�9�[�H,���h�ˍ�zR���#��O�?6��g8�v������݌�2���Cjxpq��v𚄚�d������H��b��e��Ȏ[$�
j�:S�R��\��0V��*�Y�'�rB=N� �|I�Ա��s?�~�|ے�o��l�����.��R>M,u�,o�2.�F��
d�$4���k����'�"�4���+���Z"顅C��RDL�``������k%ޮ^�A�h�����O'�$��	 	Y�:Qbo�W��X��ks
2"��_K��&��D���̥
<��D@�'p���Z�c�&��/�(=�[���i��M�PZ*
c�7����Z0�H�cR0Y��	Ⱥ���cAnW���� (���^j�`���XIӅ�� �y�w.ʝ���DhF#�&֢����T&�]$�����W	�g�����"詷�rV��J��J<��̤�(jR�Mbn&�a��|�;_� �Lb���!�@h��	\䑔��������$�>
w��z����NX:a��|ɩ
�i����	<p'�H1^�F`&6�����)X85�1�m�O[��4a�d��b��o�$��-���h��
�^b�Ҹ�4�ː;� �T.���k;@u�P��LVX߭���.%�գ�1LƐ ���]0I'7|�ϊAc�J5n��/��3�j�I�:̱��(�"P3�;^�S��q�8��WRS�S(��̌wx��Z*i�LB1�$3��h]B��mSy�����i�q��*�>1fb>�!'���Z�L� ��:�鳠�k(�dz��["��/�r�8PL�Z2�p=�D����O�UW���<�Q/P�t�������B�?NN�y��o�����~��'���OtuuEg���S��N�M�P*�Z3�pk�Y�T�n����p������kc���^�e)���yx�W$����|��n��զ�t��B����ިE��}"��Tr	�ˀc\n�^W��KzLp{lJM�MRUA� .rB�4�.Ps�x�+
(�+S��q�?�;���k�e��4�U�2�A.]f��%�O������+:9>�۳����s&z/[@�n�/��B�߿��ǟ>}������#6C㘳���^1K��U&=0H,Z�����'������wV�P�x1�Q�pi��9�x�ǔXl�� L�f�*Oz�w�63�u�p�Z�Z)6I�R(}�\����J'zNo�m��Pd@���'�A��m��dB�䣉 ��B�|'�ֈܪn�ۺ����7F��H,M�~K�u�[H*��֢�E:G�&8ބ�� �c:=9����v���*�	o�\)֝�\0��.i��܄k*����DHŦ�%�u�+���uz �1KKK��"c� ��^;��Y���aT�&�c�ƛ`��{�  8��O���C�G]�j�3ҕī�I�ZQ�Ҋ�ť���"������H�78,1�^�9$t�"���r �4�\�k�5a�耈��K�kA>f�O��e�j�NN��0�%�2����1o3_,�o��î�����a��	O�XrG�NO{��Jj�Tl�A�p$8�Ѵ�s���`�ˆ�rq>fi��z�^�)�~��;�j�lU�k�������_���}��]�������M�������g3����fK��rM���| ��( �{zqft %���u.��o7��q�O���;Q�C�g��Y0���I �f�5��Tŵ 4��JP#!
2HK�8P��D]o�x=���X[�vǹ�R?#IQ��of6[�L`��1��n�p*h����	έRB������}c�+�2���aK(\������Y
@ǃ��v)��Y�W�2�2�!HB��\�I�=-ws�Q �p|��f���W*�0��1?qf�&!W
J�b[��;^�6��$�V���b��ʢ��0�<-j	B.��R��Q�3o�S5�
�Fj�k���	�$뽷�q�	ɤҚIM���Gm�k��z�]�_��Nc>A�p��>S�z�<�Qi) Gd�ǣeZ���zg&n�g�M�pk٢�$�r\�k�c��,�H۠�LT2��Y��L΃b���w����Q1�V��zG�*��ZDqW�[O���@3k_I�4�`���	s%��aޗh ���%��_s5���nnnZ�J���-�3Ё�y��}��F߾]2)�T�����z0�TqL�e$�����R�D<���{���غ���_��1�p�#��MH9�����������#���ځJ��K���l��-k!���Z���Z����
��\*�b0g���
!?E�o��a�}j�E����fE��/8X𬕘&�cV߾]	�� b�ɭ`0���p��ӳS�X\�l^��8�٬�� ��>���޾}Ӟc��ת�w�]$���n32�Tf�j�G�1T��颃��D�A=P�sM*�4$u�"����9���`��*R�ⵒ���K�~���Ҷ2���Xe��bfP�}T�T2�f7�m�p����f��.ES�[E#"5!�A�{#D��WB��^�%@W�`5ǩ�*-[�w���# ,]��|-��Ԁ�K�G���->_�^r�D%�r��������[��-���d%; $p��#R���h���dB��3��e���Y%�u�I�,֚��_3�%����q:�HP�LpY>�@�9�Ċ��NL{i.'��4��E3�Z"|B�z$�	�`"�<̱Q��f]�t�L<���� ��� �v*�,�e����liA�/��:$��h���}��H�?��ĵ��q�����������M�惂�P�޽{Ko޼��?˥���F ��c1_3�LK:s�q��#�K��;J*�ti�}��A�I����w*�@�D���L�7��P�J�C���-�@ɣ8�v���m��j�D� �+����yx�n���z�m,,5���1���M`��^�H^i�/Dé	֕E;����:a�±8��lLRX[��aU�������%��"~���H� �SO���i�$9>gAK$r��%��H<v%�J(ӱV'>a֪J �L�ܠ�?ٽ��4V'�|{� EL��X�iCR	�\!௟�1����P����g�=;@A�مPP�hxyE&��Od��� �Lf���$����pj������ܲh�e�p 0�&��X�wZ/�� P��'�	�@����Hڣ���A�*֠��7,��f�!�� `����D$���:Qw(�.�D���(��$�{^N��5���*SZ�����I{F��70t�Q�j�|1'�UŒH6 
'�f�gs�+</��&D��q�y�3�;��PV�4���Vu�m4;:Dk8�A��r5c�a6����4���Tj'C�Z8�j��E�Nr�_��-u~ZK�r�c� V<JV�8e�x���j�N��%�����M�l��g��Z�W��5!ew9N��~�97�I��k��T���(�+fp���/�ޞ�XK�|�+  ������ŒúXj  c=�� "l�Q����=O�㒔o��� ��� �m#>("e�߂k�a����$X���H�Y���s/����h�K*�H�jT��w��`�D�:8�D�j`�g��ͬ>�����ם�z|L��s���
���s��"x���vЀ�7S���\�c���D�Y����%�[`�l-Q����V�F�X�7^lƔ�IZ�O������)r��cG�� E<{K��K�9@�#�š	�eb���H6@�d^Ui�Qyl�n��|��a�b�mbu#�7 2A�Xo�*D?G��ju�L��-�N7 (�6m��~���.faۏ4��A-9��5yG�2�Ci(��sH���
N��G\�T~2X����_а:�p1�*�p��o�Y_��j��(���#�ϊ�w�y%}� �~.�Be�f��Z���|O�L�SVi��Pr?ұ���Vdk@�L�3��m��Y7�a�­
�/ϕ��6�l
��N4����h�ɥVv܏Ha�{�U�Pt�M��S����m\E�Od���]�}��KM��1��S.�:������G��K���Ԇ|}�ť/����'�9���4���m�k�<7%�Ex�ҖS��c<Á=�usm.�@I������2s���I
$.$ o�� g�/-���f�6D��H:A;|@ٸ���D��ݶ��~�벡��9KT)�˥��5�:��s��P��/bZ�+hҫ��[$j�SI�!��+���l�YM޸���ߏO�{��KM�R� ;�=3���^�a�[z��F�I�=^�a
��&n���ɤ�p�8�u
�����v����N낾�R\t���i!ӽ�\dqB3d>�{T��9�'�J�OP��tX���5����qJi�`J�*}v�����D���t�_3{/�J>�Ǎ�b$s3�s7���%���4��� ���bP��	������l�r�~
*�3q�:�$ۑ�?T�k/�vT��A6�G���f���ӱZ��0n������\"|-���d����
��/d�uH���W�@�&�|��U�1"�e#&��*�M�d��2,=�g��gIŸ7� ����)�J8�y,X�Ss����8 �ԢȇH�d?F����4��DҠ1�mdjU���g
���r9F�Г��a ^*���D��1�RT4QGЌ��jհI����������<d����ՆL�ԑL:�P�:p(��M?�x���PZ���؍���OU�����sA��Ԇ�Z֤&��.�PҊ��`��{��bj@� s��L���~�bv�(��A�&�X��Ɯ��RnC	T�]�� �G$]�Р1K@e1��iL�u��
��X`I��� %���-�9_�d1�{o$� |U�G�;|pJK,�υ,���A�p�G��	Ɏ�-�2�������Tn%-d�q�ܻ]C��쫤}CQ
I%Sq�� �dΐ������&��ݮ#�t����6���G��,�F��P�LlN; Z�Y�-��ML�>HhfpY���B$fI�cb"�'ed'��%�ܸ=�8y�#����c��b��ӳx��c[�� �rJ��yŃ��H� �`@&l��~2�͛�I���Zh��[���
&e i�� ��&�DJκ�c���;�i�KNWE�sٞ�:��IIY�P|	P��)�$�@��aO�'X~�)��;�`�#b��~P��AJ_K�!+�"m�$�D��,5~G�O�%j
O��H*H�&#&�Fe�U��\�(����_ه�ݯ��9?,�W��*���,X��A
���S���xʻp����c^�OD��+����*��$+r� W�W�2���=��4;[E��5��[R6Ú�ɡ3
���rT��:�=��� �
d�դ�l��	�B9��
�"���$�) (��i�8�r������oE����"Hn�1�����7u�X*� f�a�Z�,�C�I;M�����kN�tq!I��8�7.czr|.:������BĢ�D+��3oU�y=>F�2�g��M��*k�l�i^n|���ojQPL�N�Z洞'�޹=;@�ul�30X����$�Aj)<� ��8���аL]T*����](�=�D0�|&#�)�z8.�EE��A�>;C��s.��@>����M'����˯�"���~i�3@]�j��E���	_��?��ׯ*54�)2V5r�ʃ����U�hn�q��(��
�I�LUO�h�r�,��}��$�VP�R,�P�H%�<y�_͏l(�� K7�Z���#�i�
��v1�;����� ly�mF����H��c��P�l�����ٯdĠ��VGd�����@~������G���_[���3����u�7�e����������?���FHiP�+�Y^�zE����_��ѿ�ۿ�6X ���B	^{n�zD��?w�[�[k�X�<ށ�U�ۋ��ϥ#i��}�7�w[�g�x.�J�����S�[ͫ���P�"�2P����uu�l��~�ɉZ�J>�$������o�/���H�1	4K(-0�e�HKK@ ����P�..^q�s��o�'�|_�l�׀�A�~d����c�Xj�E^�~K?��7������gIu;�11�,Usz䠋ʎ��;�u�l���8{��� ����>��r��s-{sk[��Aq�ɶ�����8�11PAĹM~iy�f����0�>��Yc8���,<,b���:d�j6���·ꦃ�;J�Z�Dfz�>�#K}�N͙嬖2�	I��ϟ����>M�}����`I����������<N�z����t���ꇴ�\��͸�(6/6���>�#�w:Dm��3 �Y�%��Zk�7>H5��s<�I>����q���ԅ)@�B`�mbZ䀼�1i)��e_3�"$g_sz�Zs�kN�U{=g��qs�J��	U�䌫a�%
A��0�]_�0���=?��>��p�%�͒?/�ͽv�)y�I�Cd~D����%��u�AW�b� m$jP7��a�^���p���U���͂�*�#/9K`�m��U!��j!^-Ԧ�$��K���.?J��%�&�'���!Ј�!�L�ԏo��Mz���|�|��[��D��� Y��J!�%�R��)��4'+  $�������������||,��o�ʵy�jI3�hz����޻�Z��gB���}9�̓��ꪾU����0�H��̴���c$���p?�^x�1��̈�[���-k�ѠyC36��=���ʪ��<�}�X�￬�"v�}Nf�Syv����}v�#VD����������o(�����D$�شW|~��s��ĺ?k=d�����&��	P�.-�R1��EsSXo�Rm҇/YN�y�,�H�����	�ZQ�#̙�� ��9p\ ���`8��Ke8T<�Lm87@El;��drN�A�����u$� tD}�sp����O?�E{6��'�����+xb.u�(ka�u�Bm�~ky��9o�ug7!ًnm(�}K�\�Y��%��ibk{��Z�^SP�k4�
0B/J�B��Ұz6RS�s���\�ܥ��ՠ��Lm`,�N�,G,A���� #���ݻw��':�>C�{����%�Fٔ�� P�/����� )/�f��@9H9��B�b_~e��Uɺ�W�L��"M�;�����m�H>�e[�	�����ܟV\����4 ��)o1b�@4/j�0�|��OVx^P��e�������*�X2&�H]��)�xM�m�C�J�@JBuQ����?~�8��a��}��ۦ�< ��	�G��96g>[DbZ�E�+6(  f'�'�GAmH1�'\d}��dߟ�������j�jgj��P�	�K.�F y������h"��4��\,)~�mI��<[l<5-@i���ڒA6��Ð�`J��6PV5V@lC��Z2��b��Z�쵁�Vs� ��Ljݰ���K�jj8c<��KI�zQG�%*�E�թ�p��j&+���X��B�;99	�ʣp�H����@A���q�R�~�}�,pp��x i���w���x���lN^����_7���V J�{�Ӛ�YS�T����h���6Fk��Io���2@���FA_4Mt��>��[�*��`;���L��T��$�H����s�'Ø���-D_��̮��6KN\��I� ������
\IO
	���5��w�v��r�R��<x@>`)*
~���D�{�����Ǐ���!�ޣ�ѺFn#Z���s�^�Ͻ<(��E	���|#���v@eێR�r�57��2@!J����z��Ӑl��j�����g�g����u3e#)K(�k��	�RV����Dl'��X�.���%�:eƘ�$�4�n�j���$��T"����t��]�F�=��z��٧�'x� ��Qa`ew�N�>���D����/1�M��W1Q|�V��:�V�\���@g��%h�=y�%�l�Hn�M���e��#� �#pQ*t2�F?�^�=�8�Z���]�����/Ι��VO �\���V�� m��/�R�l��q�2��^������Vs�)��\&�YCUy�?L�*�q�X���=���@MGl�Ÿ��-j㴼Ľ\�^g�����H��0��m�.x���S1Ik������5���.�)>U.�ͼ2��J�D�*}4x���+�=;��7�K5�\�KjX�|��CTu,ˁ󂓂ֶ���%H��)	�z���� 	���!��i�n:E�y�n`�����1K;w����_�i �à�Z�#k�-zt�4�g��^��ݥ'��\�R2Fst��u��g�<D]Ue���\���R��(�9xTx{Vy��,���$"b((�@A���2��b�,ۊ�Q��(�ϴqmc�VzI6b�yZ
����T��8Oɀ��F���s���!Jb[(Ѭ뾌��;���!+\�BM�m`�Ȭ������рR�4�����Z�L�=���i4*���Ћ � ��ï|��Ê������=�f���j����.5n�q�MZ��v�r_�u�K�f������$�ҜJWu&� wYZ�,���yb�4�ƛ꩹kZ"�	(i��DY ��p�R^�lE�4��(zU����Ķ��B� �F<���dH@T�2���W�\��E��)ۮ�ܐ)�I*i-����[��4�A�޼�+��s]��çh(��|]��@S[6QB3nG+�,���{�k�um@!�K�ku�KyP��\�8��O��в�'eA�9=x�lݖ\��&�'���\� �;$��
�jKR�*�(�M��Z�
�ٔ��h��>�9;��Gg����i�^�L=���zY���^!FZ^Y@��à��e����s�����6�k�+M������`�k��.x�����E��|�Y��:��m7�&}{W�[Vg�Em�������p�}��̒�ѵdC�ض��r>�0e YP�����LB+,3��\�O��Z�^����f�'Wl@�o�R��eoo����t��~�)=}�\x-�H�4Q77ԥn.�u6O�@���Wk��d�-?�I~^�"R�\<G�~y�G��$�C/�r��-�4��;WkcR�L��9�I��������� U�-%o� ���1��Pݵ�xd�\i'�0�ʫL���ڞ�)9��)} ����;;�V�8�����;<>~�8H'�lt�Ex0UT�nR�g�o�d9��r�����k2"�J@�����w�G�����%J�nm2����e+���hWZ�G͜�Ѻ��*�a��Rߘ�(��s>�ͦ ���s�����s��E�Pf��?~�kĆ�fq�Kn�<L�M�dIٲ�'�{���ϕ�T��X�ڙ��;���kމ7-���hԎ�u[������V:i���y��̔%^}��ʓ��a�xk�Fc�o�І	�LYlu}3j�Xh��5'RB
���}���s�L'���{��>�faS��׾F�1�I]��z���xx�-��d`��=��䭭��9R��>)�����gI׍�[�r&�����g��0	��>�6BN���EX� E�d��<S��yZwW0�ww���.�G�N�(�Z>���s�Z|fS��n��O�h�|��7�/��9u�E�p���t]��+{u��?��Yi4���o��Dڂ�Vy����F#:=;��m ��+Tǌi�k�}��O�T�����ۻ���l�+����Ɂd��V�"��[_nƪ����:�I��K��󚻀[�u�۪`[2���	�1�2���܀�J��̆��Ɏ�?p1 (��ݣ�)<H� ����C��Cr)��5��y=@qk�_�=�����`��P�9����`Ş��D��s%H	���6��Zo[�q8�O�M2�ʈ�`���ȵ��[H��ـҳRـ����(����?K�غIߑ�!�h�*���W>J����S���K�I��`�$�!����-h�`�nb��qO, �&�Z^����G�Պ�^�ޗ�����y��,_Eǖ�Ͷ�`"�����<x��LW�p�S��&����fFY��PjM���&'Vr��|���uJ�XO7cE��xy dpNڅ�WE� �f�#��/_П��ص|�yhq/�D}�A�sR����!%c�z�*�H�>u�҂���]��8�eE���m�4lm��j���fx�nJ�X@1�q��-tj3�z�|V���4�`��w&�$���y��Qܥ|�9sRFa��b
�8�5]����@��~͖���#�3XX��I9����yܔP��-��ˎ�C��r���n���Jĸ�X���.)e{��鶍�>�r`�����i�`���S����i�H�X$������H)n���8����S�f��ll��ۧ�M��4�۔���P8��U���g+λ
L>��a����j�3�����>u�� I��]�ȉu��XQ7I$�z,I�������6P��`}��s�+g�r�P�J(V�K8��cżO.��+ �š -�N�t�t�H]�hV�/�x⠘: ��k='y���#�^IkI(X��Z��&�yt�|(޷�+�I�������N��n��ܮ���K�e������~6PV6�cfɫ�C����1��0$��T�|&��G�k����e������j.�~x�"�����hzǩd�׉�$��X�J�ƻ������]t�v��Xd�L��O���ĸnru�~�l,]��.��&���3�����yu?�+'i��u6Ef��΂KPӖ�^{j�\�r����>����#A��1���e�Y�`Y`9�H�v�xd�����^`��<>[�s	@{�yo���|3/H�����=��3�"��<�˨�8�2d����5�1�e͊�'��M�x䗮�ۦ��k��ǀ��qm)+���C��i8�⥍)�a ��3��wV�_��Z�붮�>~1�P>8\��!*K���s��6i,��mӠڦ��]��W�B_������&�Ju�ww��e|�����S.�uvv"<�f��!e~jB�U�~v�;��k��j`�$�ݺ�6�9�@f�;]��9gp�ڑ9��4yO}d��1�=��ɄG1h�>C>X�Py�a?"�(�iV�h<�WP����b�� \�������m�6�ڙԚ��x����>1hn�Ym)l�eÛ>_h�Xv!:�e��a�9ڀ©K�$�dԛR��Zsp�78�I,M����a�;�;��R��K_�}���}��ߥ�O���	�g���m)GǇ��	��>}�I�Ṓ����Z��匳.��]�O/�E�&�c������*�Q�,�<Q6�R�j$�럣9��X�d��`��Ԃ� �v��j�E0'T�UKz��KW�h�V+$��oDc7����[F�v���#Ku5�I�ѭfg;��ʐp���a�b� �ŕ<)�t &M8|G0Ih�╩��� )�����%�D�q�J8|`0�(� &w��a z��{t8�u�HTHk0e5���3�`�`_�L>���A�{���q|������$A��P�E�[<�
+o%�H���^�#`��{����4IB�Mn��x�E��&�}$�L_�$��]Jbu�l�)$����
�+��m��@F,l(��{�n �9��99=&�(�P����y�v�����i���	{W�N.R}������I�޸%�J R�L�62��,��P��жd�@P�H@����[�V-\��MbH%�l�eI�5H��(��.�>��p���ˠŬ�1���4�d�3
��@��ϐ���9�����i��1�D�ߥ���X�x��S��|��A���#�'Oj:�2C�ҙdkCy�Հ4�����o��^���>Ӷ h�nDf�b�iT�s+>k]�:���eϓ�ґ����^�O��-����Uy6�m$�ĶBT�uq�8,���}0��d��D0w���HZU�s���I�-.o�Y���Nr%��K�����za�"K��}|2��T���{��;�0y�C�{��Q���OX��C��]���6&"��q}� $xE�d����خk�2��ի#}�IKR�y��;uœ-�U�33�7��79�\�����ڠ���b+���K�I|�=�B��@Ik�X�k��QE''[�;��"C�b?$��o\��i��ٸp������PP����9��Q� ��w�M�R���(�ԍ~�&�,Qp���̊=>~��ģ�{Qr�r��\N2���E��V�����{��~�s���M;�8��	���w�����ץ���}x�fʊg�F�l�Y1'���u^Ĳ�%*yQ�M ��� �G16F0IjŦI���G��	�
�17#�!B����.]a;99>�ݽ;��/}�@PhiҒ�(�D�sr6�s��u.�g�>�GD?~D��s&�H5j[S�x�
�bf�^�fr9;�eZ+ӽmo`N���g��Dlm��a�L��h(d���~=��=�J�r�>.Uʮ�O~V���OAJ�,i:��Rn��xʟ�=D��T�ƌ8�e;�����p�5�6�F��{�^.Kj W7�r����wa�O͞pL�&���ARy@�]�%�t�h�1��GɤPV��e֫��K'��b��Y�e��fm�[׌�9#F�&�2f%�R~�$���>���������9Ncz{m(}C�DeV]ª?+�{�Rr�MȿW�>@ ���H8;;3���P�O��`P"g�Rm@p��ׂ�~Po�݁{�נ�@�
cw �7��^O�P��d� u�y^�����U�aSIFX)J�zy'�έ��t��,�>U\e�O�_2��!�2���`�=�y��_ӳ�$�s�^�m4���I���p�yy��n2���RHRVf�%yN�9�� 1���}VS����L���;�x<��# ")�^��ξ�<��xEdPr�O�6pV���nH&`n��P���p!//�E���9{�dE��L.+]\��s�3\�Z�RC.���P����u�}%�&�NN���rm��s+G =@¿���J��w�S��i#,�(}��^���
�5�����;�y4��C����J��D،�^ɀ� L�IP_l��3����z$�/G�C�D���D�,mL��{�w�Ϟ=���������p܅A�j�h:d���kϟ��期����0��i�&��1�\��b7f\��Fx�컊�4�m.J��"ϣ��m�1+����͎��q:�i(��I(�jS��� $s���9�E�B9$>��ZC��J,�4bg �{�l*A
A�����DH"R�NON�OpC�AL���`H���o^���,�����c,�k�5�iQOբ�dE"�;V���׼�V�Y�ի��g���\n��A��۱�����s��>��P�r)/?���8�P|t?���6վ{�(	p�D(�V�R�8\N�d��q��$���kƳM�('*j*5  ��IDAT�~���H F`���ЂY���Xt3�@�6�Ċ��LN���qE/Xr��&����Rڌk!�dB��� T80P��7����4v�p�2l"�[j�4����)�KFʞ����$\���BIJ�ծ�4��e�E��p���l�%e��MV�3iA:�� $�| �)#PKi �<��&�D���A��b��*�l:��a'Y,���D\�3�LNNN�.���nb��ש�#q'��$r|�΂Z�%=��3��@�J^ٌ�[qjK�Y&���o ���f\���r@�N��E���yOy/��m*��U�*2��JL� �fJ<���y�cC[�*^�(9r���b  i��.@�{#���(o���82�@>��1=y�$|������=��ix=b[	h�����"�uU:װ;
Y��?��$��l���+yi��;�w�
&Ҫ՚�4ޣ�i+�+?�e��c��5ʚ���!���T�s6Z��e��J���>���S�]I����^y�=i��o�ڳ�����K�h�X犈KrJ)���a�Z�� 
������P \X��
����Hm@	�����:���~�s8�<Ӟ?{^�{b9K,�tzF��yP�F���F>�w���^,ʠ^MY��\��H*՘>��V�֮��s�� $��\��W�PZ�ds@YJ��殈ѿ�cɡ,����]�[�u��msE�Mf�K:� ���-%{x\�a.��=	��ɭ�񶙃�1@R�*X���vu�)Ol(�A�L�8b)�<P= E Z����'4���kQ6l�}��0|vL��i ��N�@�P��`��K'|�5*a�l;l�����1�Q�܇V�[#��y���n��Kz�!�\�ylT����E1wl���3գ��O�ض���O[B�p�B�ͦ�r*�E��Y^3ǾELGa*0�x�{��F�;3(��m�c3�+����Lx�4w���Y|,nmj���(�*+Ik3��S��G�f���KR��k�X�+�g_2WLT��4L|�`���]D��vX�$��~�L��J3?�O�L�|,��bYp��Z&�'�'�.�|\���I�ܸ��WeR��'��܌���h�ҠD�����)��ْl�"���H�/_[�7�T͕/-�v킗ydx����������5��(�����ǿ�on�S� �&l���eJ�n�fc�>�L��"�%��J\�r"S��T�mt0Q�Uu�����TφOL~�Pn4#��q�����X�y*v��V�\W�㓏nȓ�ZIj�ڝ�5�W���wH�Ah�� ��bT,!%{�dV�AU�@��@^A��p'�Q���%��6ȻL"�F��&t�<�t������(zC��bQ;�ѷ$���Ԣ�j.�A;���Bqj�k�s�\�l��Ӣ-�Pa�ɲ�b�o�Q�nm(��ܺO� �XX�~Z	<��+pi
I|O"�����uZi��$���1���Ҡ��ʂQ0����I-�� AjE� N�Ll4�L&[�`d�D���� ]�� �u����Q�&�zG�g=zeN�4ET1.c,y�5����A��ݓ�9Ot�M��
~!�E*�ӵ������޲vmD�X@Yo�k��.%:�}�9� 1�9_�T0�ud?�&���"��H휝�bi,Qt��T��l� �2��+�[��n��s���*�&_�����d�4�{����ν��R���ݦ�e�%ν|]IJ*����G�#?�$Z���s�5�Nd�en���6]~�"���7�m,��[�$2�J���ME6��s���Cs#K#��@̌����4z�k5?S�陻�l�E�������:~� �Uj9���B�sxn8C���*6li0K5"�QZ�^E)c�vW�˘O��� /FK��V���~E鳧��a[n���$�µ��V0ݞ�HY��&I���L�����f&h�(�����f��{_�m���D5f�%
�yb�ٚ�$O`��I�v�.�d83�eZ�p$"�����4���y�Wb�+�h4��HU�� �ՇI؇�ٌUq��J�?9W�kO`z��_��ܺ��E,M�:��E�C��ז��$���lp���;#:Jh�v��7K�E+%�\����Z�$n�����_���v(�E�[r���2�#���Kl��ǒ`ɲٛ����a�`A���\6�Z���nW���#�/KS?�x�������e�H��Db�����4�{����Z7�&�a�]�N��OJ!׏~/w6Zu�(�D�D���b�Hׅ
�R�dbǎ�G�����-�|VmY[P�Z��ą�����Z{U[�%k�t��"MT&�f'i4��+Dŧ���w[[�_�S��ec�S�V�1F�L�w`2�v_WHX��q�h́�ʊp0Ԣ:i�,��ižU��Ռo�I&e�/�a�v��� @���-�В���*IA�6�ET���;����6��?}w->��mv=���@��o�(^8˜5�R�}Lݮ����l�ל���-�G�vB�H|���,c�%)%}b6����� �%KΡ\�cې���I]]V��y�W7T6g�).ob3�'�5.�ٹ�f�V���K# 3".��@���sDzf����-�0A�X@���l�32�@WR�[QƁùM����`�Y9��:+$h�+��E�(�}(�~��y1"(ȑ�H*�A�1�R�l�&��^|ަ��Φ\��n(�u�߯�;��W�r�g�JVe_��ẆY����oT!)����򱋊�c�M���<}��U�<���^���L�X@��@$��1�C'�W����AGq�H�'����xNY�-�b����]X���آ�S6ٟK�.�ɛE�b���ň+����uռ��C�w�8�SO������>����r��{�����4�����t�����w{T������ZQ�/,htY�h�բ�����e�N5ȷ�q�����a�����<�@���n}��=d� ��v��B�����6m���C��lp%,���"M��_�F���Qu�(Rm�&W��,K�~iF���&p0!���U\P���}z��w�����D��>y*�Z�e/�T����?��e�¾��B���&�t~��m׍�=~w������W^�6vo��UZWf	�|@}�7�m,�D)d�9�Ē,�b�� ����q=�����;F��%f�&��&���k����W2Ck���ܙ�����Ir�Vi+�Id���Gq��(�M� �9ýG���ݻD/H����%񿷏�����m=�Mz�Fs��M}�h�"-�u��A>����t��U�*�J�����~�-��}��P�\3IC<+?����4���M�ٽʅ�A����,nN'���7���b����6� &0�����^�=��G��h� ���<�[��߁���;w��@�������� �"�q�w�у�9	�Zɰ_QX��*Gs��s�*Ͽ��w}&�y��ȩ��i�P�&Gf˱�g�ie�D7�X��j��5K��P�T��-�8Z���/I�7�*!�_+��ȴ&O.5Ժς�\t	�Y]Oo:Z��%�h?)�{�'�#�����m��e��v0���=��� ��8�-*�����d�,[s[Zgz�[��r$���m�tb�E	3��t��A�0'����细��(����ieJ_�J`�I�}�{�<��sD�p��-���&�I<͢h!��!�XB�XOE�X`�A664�f���3:=;��B��Y������r9N�'(yb�&��L��a����)�!��x�K��?ǃ�����0 �{�� ��N���T&�zn83ܧ�~�i%��s�+���W��M|ݳ��Ьr`(fĵ�t"iR3�7�D�W�4� x(��g�Z�8���K�Y��"��\�,�C�@N�z(�qzzʒl�2m��vn�S�������|ie5O�����d��CL�w��b� �l0٣����ּ��wikk� �����B�7��D:J䡕���&w�yl�����&K^���Z����sOG����D�j��L�.p�G�D�̾��-��c�m\Ē��m��zAKޞFKl���C�G�)�.�(�� #!a4$�Y��&1pCg���N���S�)i�0���
x�~Ξ$�A�	r,�87���`+�Qgy�jݼ,�W������5��Z=;�������!�k�Q̀����w��sp ��;�;����̜3�/K)�W"��k�ܠj-�D͕�R U�zi�ϟw�n��a�ڔ1�H�~�=�	� ;��h(="<Kw�̜D��o��B�,��;�Y�uٷN!�%<�^6�m1Z���Lo嚛�LL�����d�O��㚆������/���A`�>� (�� 챴!i����h�^������}Y���s&�Zl.^(�U�E���5��9�ۈ*�����ܥ�?�z�s�h������ ��^D��������=���,$�l���i����u���d�b_}��Vw�:U_�F�4���B$�G2Y�	��v0�o<����쭨Z�Oyl@I�{��(cǊ����&�i P$�\!F{����&N)����l��~)�m��^�eMo%�7��N\\�P����B)i���A��!	5�(@�߿��d"*��{��M�B����dS+m�QQi�t��loѝ��rLF��s������_�w��\8眫R�)��V�<�0D��H[�Q{t�����)���W��Mں�f�&����5��>3���u���u���O���㢴��^R�yՆ�sB�0Xf���f6��4�b�H'K(��9����<�
^�v��1��k̆�B�>�T���In���9(d�.�b�+Ճ#R���^Pk�1(�=l#;ۻ���_���Uz��w���'���x-&@� +? �,���� r|rD����o���� �m�<�>�e���_ˌ2@��t�#�(�kmQ�
�3�n����֜��l�	/EA����j��D��э�ύ�-�jEЭ�%0��b0�\d��8*U���BEj�$�#e�.ŕ]�%���j���p���llE���V|З��C�O�<�g�E,G>��|@�H((�1��ET:���c.�Q�8X��ӱ��r����e�LRX�R߻����@%�ʊ����ͅ�$K��~�'���㤣�Q��q|�zw,�-��4M�d��%���:��d�e��������7���_���}ڀ���Ҷ�����51�#H��At��Qǆ�̌~2�E�,�
L�PFj�`��|!#�_�xr��x��~远9?7z1�[A�c@���>`��?����'<X(�����3zqt8��[�c���L�b`�U�r��ʉV<b722�5Lh�(�uؾ{MWؼ< J����DtK�5Wy�IY�[@��h�ե��Z6��e��F��x�����1�)������nU��o}bj��Sr��X+Ԡ���d�iQ��J?����(+]��='����@�T�(����������*��4H.��Y�7*��;��Q1�z�N���6�θ�����6�m���y+��d&I�8���2s6f�� ΏHX�0=	 ��9�*��
0Y�%J�1y|h��zI�u�ʤ {��!r)�2�g����Q[Z�SiRٔ�'Sg�i���>g���&�B���j���׆~���"@p#�y6P�Z|�bA%N}o��2Hk�zeƬ�B��~��X�¥=k�R&�X��(���R��&5	&�ӧO9SL+3�Е��8 ���p%A�c`t����}��W�GѣG��1w9.�����T 8��N�tz&eR����;�Z# �`�3��}S7qy����n�l��3j{�z���B�D�����-{�����%����\a��A�o%��l��ڱ���e��#�К����@�z�Ra@�V�ϓ��\�\���+W�񴮱_���#vf+lp/#���>��7���ײ���u4W."�79/��\W0�V�xƩNNOX��ʄ�8��x�R�Ŝm'��Ny�&��Տ�j���f��m��͕낛�4|���ϳ��U���,D^��RR7��]m.U����KS�J�<?���m�T��%^�x�$@p7\�	�������B&�����UJ�⡋�SxGR�/e2���A%L���� L����R�;�р��|؃I���$���py��8-%��~�$}��x�� Y���� EHV��b`��S)�~z~���-Ut��0 
�2Ҭ��:�q����L.XH�}m�j��HY�ցH�����̛���,+��ķ��%�Č�T�5�/,Wy:�0}��ߪ<�����탌>���O��qN3�[�*D#���Dk-�5�`� 'd `3���%L(V$ y�
������|,���+c�B~R�)�s L!�N�8T��G+C:9 ������Gl��(PN�� Bj��T��v9�>��r�f���Bi�'aw>]��������&�j�eTۛ�,%XcۙF�����'�U"�;��GZݖ��'�d�1�T3���ɻ3��mc�]�	�Q�,���7����h�֤Z�P/J��% 6L��h�c@R xL6���x$;�zF0��8l"h�r0Hὁ'����$�S�Lɇ4���0�:G�t��TG�&@�*���W��p	K���/�в��3�T\���=/Ԟ����jNs�iKLt��$'�u��l��+�$��@$w��k�ڈݦ:��[�u6�.�NR��$��L���5�|"(Py�;M]ɾ���	$�> YTJ���J��[��6H'w�ޅˏ�y>H �jb�ILdX����br� $%�����8|�����<zi��G�B�⒥$�$:b��GP�V�ɘ�(D�޹4#����7��������>�GAi�_eKh�&j��'�%_�ӹ��&&n��]oZ������t��Ƚ,"?��+�P:c�B	�ɂ�t�t���,[wŕ����ȋtY]�q7�^
����t�nX�����찑��c8R�c��%�6� ���$�uA�kv�H��wX��?�#���z��ӏ`8���\����bd�ͥ$��� U���V������"��>	�")�u��m��Ӓa]��z�wtt��u�v�i������J-L�1���@�*Z���Ƴv��Moo	��-��i�m%�JR/%�c�aI���]hd���}�_�lAi(�D�Z&�ӕE4��w�]A�v�kDꁏ>���� ���_�}�>}�ꎬ�5��x�D��l���^�t����hyB
&z!�ue��{�oH��(m�\B�~H&��%�<�8�O:�T�u2�K��V�����=J��X*���,����͐M��9@P3�� ���T����RmU}�(ߖnLd�Q�UB�5�^{[�6���dE���E�F�aɤ�:Y�mU��m؀�w�����Pj$���5D�oM`Y��'��������#"���IA��%�bPq*&k̝c��Z0`���$��]��\�r ���8!#���D�Y�I/8�ULOϐ����$��ny(�ے���?ׇ�#Y=IJ� &�"���he�j�U�MX`��'Pï��������
/l'M��:�A!`72�E5�x��X���%�Т� Yh�HRi|N	�]+W��X*2]{��*%�x{2�l�T5Ī����fCWrX���[���{=>mǪ��)���9�w�R��:�?x�x���Ƌ�[�?ѫ�XY�(H(S��m��k��P�Nl^�S�4D��1�%%_��mjم,����$!U {��0��w �|�0�$� �B�U�jpn4��1��y���3i��䄥��Lk*7��(,Ns�Tt�ǹQ���$/��B��E�y�fS,G�5����A�eh��A���{g��N�Mm��������1��bg�����>;O�yKL[�Fqc�b�`8@�x+P�X�@��S�]��b�A�d�6���{Y
�c��؄13�2~7{�VB��&��$��b���� ������{���dYdp���0��^"��3I�P��9� 8%���Y��j@�� 9U$HD3vSw�d@���e�t�����}��'������~㚦��5$$���+¶$c*uWJ��ړ��ϝ&��vˣ�}���u�[���eYT��E8�Z���,e��^��8,Z/�H�]��%]Yˎ%Y�J��b��'�6��xK�t��̥lڷ._@O�X8s���:��*�L�ɕ��� ��m,��U�Og���3#3�Ii�\x�ET�X�Q�	dl	���f�^���L^��^���Hw��DDt��33�ڪWB|�qAϯ�l%� ��
5Kr���q8L�^�(^�W��qotB)�oS�lj��PhIAx�h~} ZG����$r^�X�1@1Wp2֦�t�f�kV`�ϟyu��^�lm�^���W��y߹�&�ķ�?@*�y1��R+_�B/7T6PV7e9���`��R�WV��i,�KVJ�$�+�j0�{L��<�ʐs�X̆�0�!���� �w�� ��y�+JN����7�E��Ex��Xz��\$��� p��u�_��E>�4�FZ�����\�f+�W��^���ˌ��oR���}? ǻi�Y�����0aI�6���6o�Xw`��c%%��b�9ŇHN�Z�!�߀%k�|ƌ4/ l 0�J�BM'""C� �Mg��f/5��2�$���=�V��7� ?^�E= !%A�͇�J*>ƃ���K5� �v�T.2�^����l댦��%%{5�$[R�`+<N�{�T+�Q,�z;tǀ�]On����)$�`�"� ��[	���(~�}�9��R��D2��2I�&�L��� }Μ(� ��1"�xzfQ�p^fq�*���X$!LVJ�:��x1c����9�3�<�hB�H��w��Z[6^�]�Ȉm��I���{ƻJ^]�XK������R�Uqy�.
ɧ#K� ���C��JN%_�zW�lu4��U-3�^�!�6@J�l,~	ރ|�	'm�L6@)9=#8%��	�b�Q���3S�+�T/�O���-�00�!p��'�$��^�r��"������urd��?�YP]	��s(�Rr9�����Տ�Ә�n��`�=W��oF)h�Q3:ߺ�O?Ǧc7j�^<����x�S��5��^k�'�Af�`dD�b`�h�0�ͥ�		�S@�F�2AE�lj �a�N±�؈&�2���x<SWd͹Q�qEJ>�`�%�͐F�w�y�� �-R<>���?N����E�*i�:�������`�hl�9Jn��P.ei]KʇҒ|ܲ4��l���L�FT_�$!z�N���ò�s�f0��mF�X@I�[�j�(�r�C�@>	�P�s�'9�s,��`�0�k�χl,E�<*PS�Bn"2 
4�-8g
���@������	 �,�T��P����IP���=<<"Y�(b+���U<ށ�BH�N�u��z�N��p�S�����v�>�m�q����$KY�3	�U��,^I��,`�-{QKd�4I�}׎EN���������ʫk/G.����i�����֕�ͼ %51 ̤t�i�ܬ֔��7#j�jGҹp �M,�o!U�̾1`iȃt:-8����T/ �~�8!������	I
�b�V����ϔ�,[w�ކ��I<��~g�R�K�5���]��X�q�rU�iJ��<�׼�<~Pcj~N7L�6PV5.��5��K�X�J&�ѐ%L` MJI@:�'� `pzv���� )癱E|�S�1��R���h@��6��-���ɳT���@<�:ʥ�o$5�B�Gj�l�R�^%_�K����� E�CPhPV���p� 
W�m*W�����]��6B��l@�	P�L썴jA-�0T�Z����ѕB�f�bo�^lu��&�4Z(��Oo[��1�)���f��,�L�b�0�JXr�')k�\� T��X�\�o0��I�[ OV�	'kB8��\�ߛ*�س��Z;�J��'K'���ѦЋް��.�,GS��&��ʆ�i��Q��h-�6�\�1H.�%5�<Y��	I�`)��pBo��b#�,�X���7�2�I��U 8�����M�`1��m��:�$]X�j��Nu_�r��a�CIcp���6�8��4��bIW��+.b��[c�����'ǜFR ���x=::fi�:i}���E�+��|ƭ�_yYi*��
�Q8j�$"�\�_��hS�y�k¢B�)7P� �2ޣE��W�201@A��ź#��ǁ���8 ��b�o<��pQ��8#'Qr�Jr"6�$!��3�Wՙz�J�\O;-�>$�R\�8�pi߽7wņB�N����*GG&���˂CW�z�֖N.����`}1!��G�L-��1ۚs-U0��ݺ)݌�Q��M�*?V���7ҒTҕP"���|��\ks=�%���Us��`ɣ��fi4D|Κ6�
k�+�G	E�5�%�-�~/+ ���_�\�d��cr��Kd��X��TjS����.moɣ� �|pp��ܰ��z8?i��G����Yb��_u�]1)eSZLV~KA�Q�آ
w��>�I ��W�-�R��@x��J��n듞������6P�ګ��LF>_K�]����b���$[�T����I�7K�8vπd�\S��=E�"Y�(�V��Gl-�=:�z����H��)'f�� g�H]bL.���Ç��!�2}�`i���n��ϥvi�U��t�jK ��iw=�����,1%���(,A*Y���w�K�[�SNwXC��B}Hʜ6�m4��j�������id��	@�$Qe�1�������`�yf����.����R�]-�!󕫈C�pWU��.5͒��)�����޽�����/O��1T��z�}3�� �|��l�}��c64�ܖR֩.7Orɍ�iK���)"��F��
*+J�����,�+0�k��2^����V��VB�,�Ib�h����֍����#��d/�ꯒ i��2uI�
遹����<����D8�cǈk�{��n��7d��]�=�dH'�'B��B:��-P<g�1�4p��P{`��cu���������e�`�)��<6��>_��-� ���=M���/���{~n��A���񵪇)v�6.{�&A�7����D�/��'++R��������w~�nz�X@iؽ+�-Z�l[�A��Rl�Q͒昚��|�G5A �2��X]jl��`s�o���[i?��'�Wcm���@6!���$<�ً�4��,�<y��5R����O9[����g�R����ٓ���`��8�j2vY�]���1�Ů�9�r���� �k�����Z����d��H��ۣ�\�r)�=jb	�<-��\�"�f��]��Q�6m�rd9p$��_�w:�Yq� �����"E4wj���A�iK)�]�m�;�Lㄵt|�(���!"u�F�
e�N:o�I[4p��Ưl�G�h�?�3�4���o 486�M�x5(M*9S�8�Q\��Y,Q���%o�����*��=Tn?`[C��qD�Y�90��U�+*5%EVOG���7_X.j��`{Z,AB1+�s)*�*���V2�J�����,��ۗ4�R�9Ƈ~e�6�m*�p[�B��${����I#S����3`׷>�F>B.�|����w��v�>��wQ<�|��6��r$�H�V;,����%�^>��]�.�P�УC������|���q��iH}�D���l�Yڮ�E��j(��K�%�c��a�ht1�{���L���` �ɷv���������+c6y������}��s�j !�h�yS�]Ӱ� 
��"e��ҵ����L��z�Y2ck�����}K*���AT�⥵��v.۷�{%럩a�%&��f���Ԗ>�jp֍���S���2�u���ʪf|�px�+�zx��M=P�j��a��^�_j=!�-^����>�t;�̔'�0#�ʧ�~ʞ���Sum���sSZ�L�m�q>�}\jwQr=҇�ZĮb��$��s�%�6�'�-���� j�8�x����# Y���o�3qUe[�J���e*@5@s>A�I�QPsf�3�;���$���'����3�� |,]�r��~���k���>�"bn��E�1�V���m�ɤ��}$o�(K2�y.�b��H[eQ�Wx��ݗ��6PV�܇_����Jl�S��"R��x�{z�uj-s�L.�!W��^�F�jC�9:z.��	ɭ��pY�����P��Y7�Z[|V޷�����'��~���� y����5�+o�_8��Q�*�!=7���V��)A;ʶ�5��\���#�ms�����e�Z�oFXJ���9!�MՕLĀb�ںC�^fM�^�Uͭ���+���Q�F�#�2 .B��䘠����yVp͒�R�rC����7���'�K=�8���r��x��!1�̪	/��
r������O�o�T���������3Yl"�vsGP�랁�:��������U����pE�gb���3��&�W�z=3�D��rSk')}Ju %��@{Q���2����x&9�Di�>�n�#���H�)A���τ�je�떳bM:L[�[�w���^I�wT12Ɍ6�m,���4^���/L�_�cUASsZ�4�~*��H�6��0/�Q��/��4R���e\��'6��b�0��C�y�g(�#�Sy����mI��z�{J�-ya�ZJVA-��g��+e�/n�(m(QΒk��]���2��Q����5�V�I$�6P"�i��,�Q�(]�gZ�8ѫW��k�5�,	Qt��%��+LF�&<���4fP�uk��&��x�k*l8y�/I�������R�~����ev��vm�<]/�}��%iD�O//���X"�eɦ���ƌ���,���+������m���Za��,W<t����F����8��ÂO�C���tU�j��uF�c�nʆ_�kR&/l+\�������ɸ+�m�>���'�הX:?�%��S'	c%�e�"*�=��C��;��}E�F	'Oo��% �{Mƺ�ra^Ͱ���FʪV8-*�Y�]���e%aNLС����\�Q�
P���]�H�A������P2A\aj���"\2V�����.�ǫr_����
�sm*��ύ��O�u��%�ˀ���<ȯ{d,�n8ƒw&'����Kl��������`�#�d�Az�L���<j��ʋ�����æ2(	l)2�9Z$q ��_�)���:ʒ�+��<]
���<t�j�t�:�YD5�w#v�@2C����\��'@a���.IS�M�~�M�zo@S+�(NDZ���
��X���>��ۗ�����3��Vjy�6b�̮C	Mڊ%�_Sh�kޭ�or[��T:�À���mJڜڳ��"^<�"YZ�N˹)h�R;M|�c�k�f6ϓ�L~3=o��1�XQ��M�'ߺ�NK���;��6��n]w\j20,%_]��%�칼�7c+� �@y���K)�Q
xxXNG���ٷ׹7-}ʤ#s�N�1�X��~�د�W	�x��dKT7Y���}������"��
��˒�P�7�2��{�o �b	\��]#��n(�Z�n�`�Z�Z@����&=@�����D�z��&ZW���B��/�R��_����$WY��17I��F�����������]w��. ��E�U����4�Y���MJ,�Jm�:Z���7�FEV4�}\ˆTj�M�\���,���Г�-f�n~�>'��]�,�bl�V�����(��'����=�{��0c2R֭�~{Q]���o�^c�扉x��p)lX�9�f��"\�"�}Q�u��cN!��ѨD�d:F|��u�u��Rp�� G�+-�WP�o�h3d�C���^5�$�B�@�c��f�I�ű�����:�C2�T�V��I��O��h��-�7�m,���JŚL��׈}uu,�E�� |X�m�#��vd/"n�N�;r-��¶z��S`�La�|�W�t=~�c�:��w.&�it��$������ϧ,m�/9"2����dœ��0�����
)
?%�����k���]K��xb+H5��'q� 4pn|j� ʌ�'.Z7#|T{�4��o���W��k]P8�#��g��U�p8ڢ[@�����P��HD�4�x��۟fMܤ��k�uת4w���
��eGc�ބ���u&=�Z�\4&	,�OG^׳�����Id�I���ލg~M��ԗ�{ߵ*�v�G����ˌ��i.^yy��p�̠˟Y,�Iҍ�f�d�U˨�q��q� �@BQ+���Mn�\�ɰUwh֍��H(�ϷeY�}���>����մ��v�����d��&���g�j��o��2ds)�*���S������
i`�$�i؂om���H$F�:ƒ�:$���K�xq+}2��b$�_��;3DW��$��6P����h�A��V)%������u����_�Wŭx� %�%���yj���z �%���bL�Vo�ZSɝ�5��@�5�!��w��^�e*�Hu\D���l3�h��.@<Ɗ�ז��e:Z��:�$9o�m�MUPn�ڳ��[n�������*	�b0�{�n[_����  ��9��b�f��^ˢ�ə�8L�\̈"b���3�*�Wg�Mt05FX�0}����b�oH���̖������M���ѫ�7�-]�O�aJc�����[�5��51��J�zx��`���ԗל$�Mʠu�-��̡c�$qIډ���QB)(�4�5NF�����s���m�Ike�
�glF�q�v���.�x�6$�ɫ�Ģ���*�A�6��#�IϜ���ٕH鴒dk���X��|�=ʍ|�(�����!4�ضP�k͆�n%��okM��&�T�@2�%��=���,����I"��4�VJjl�cӰ�)J���F��^dD1��Ǐ����2繜ś�)+�<�\N6^�7�&��<�ܘ����H��#\oX�T@���L��sI	%ڎe�+�\0moӍ^D^�ٕu'k�tҒPH�"zou�"'K(�I�H�=�-duoH�� ����Jؿd�^[�����̛�ye�D7&��GG�!��QWe$?b�K�.��*�������4f�/ �Q(�q)�6��a��	�G$�rcAeť?�=<�b#VJ��xo%�K���O{FEV��@���I}h@p�S�$�ʙD�r�4m@I�A����M�.D����h���9$�)��e��-ڍz
���=uIB��49����F��4�L醶M���}�Z����y�b�^�'�"WK(��􌎷Y*Y��f���'5C�s��&�555�
(�����r����T&2\���e鍍��(2��=jU �Ҷ�`3�+�ä�J E�#K�RU��z�������d�M�������_��O������k���жI��r����m{C-��h�݂J/S�H-��jJ*�+S~��-xiQh+5/�pe�&�Q�C��D)�j��x,נ�$�a�%��R�-H��t2�/���>���>�	���V���I��߶�im{,�Z�8S�H�KnL�B�ݷ���h�,�KH�>n3�R[%��!�;���Mb;�����ƣ1������,j�Q'A��q��f��H⮭���`�=;;�`2��6P�9KΓ�u�\�E�^_�,[�W�ζm�n�l7ٶ6۶m�mv�m�f�V�������o����>��}ϙ��F	���-�8� rs�pg<S����o�*5W�=��N��@�k�<�!z�j]�Cɲ�&��	�@�ʍ���ׇT��� uȪs�1=���#~���2�V87S/03��}=&1����✍ρ�s�v���G`e��i~6�o輭�9^����l����C4�[-�PY��Z��,9 -�Sg�� ��ǔ�XI�J�WkWd���J�
*t�m)e)�6X��f����i$��w���N�g�d�ƪ�T�։����
����},��t	�.��EZ�	��z�(̩Z�т��i�p�^7$����W�]M���i�ݺ#�=d��<c
XY A�vw�~;Wc2��U�Vl��D?ZRq�׬���Q$�"����8|��up8"��`��)� ��b���PH���}���}�J��YV������>c@��姩���{����fLu��ǵ��ڨ��N�[�����������.G�������,E�2�X�N9�K�r��w�My�Wup�hQ_p:cH��'���H�/��w�:璪��/�Yq�s�1�T�Y����q�j�2�<E��C�!�4�2��qr�v��}~ny��uM��#Gm��ool�%;s6�u��{��Q�̜���Ǥ~3��ё�`z����[�!��e�ل㫎%��p%aH4�����:I�-�@���UY-ߜ���/�g��k�vp�I��I�BK���42b?���'27ŵ&�R6���xX�q �����l�}�|�:)�*e8
5�܍�e��z"�~.�i��H��J�����k�~5�lw��ücǴ5��1���=�� �V����{�r~��	]l����_�8������T8��YQv�n�]B����f�80��C���>�W2gKK�z��eX�I�vJ�Ů���L:g2�TV��MNi�vv~��/C���ݗ���WWA�����y6aӁE�x',�z���h�U�6��w�FU՚<�h�KMc�hm��|_�|f>J;��I�0����N��R؟ ۏ�cЦ`��^�\ ��/��Äz��=���$�
^)�V�[��A"'�伴�^����quv}�j2qK=Km�����6�?¶�v��d
\	�[�}$���M8o���b7�uQ ƃ�����7����t�"�W2���d���yU�&�V
�ɰ�e�6:��,3q�����:�����ײ&*�F�4*�#�2�+Ͳ��=N��ƞV��M�� �_���æ���LV����"�	���R��BI��L~O��޷�dw����;�!�1R�{�Mv�����cp�n�i\��I�5��6����o�m��N�`v��y�Y���|��}z��|���0U�*	L��`���tUqIr�P%\�����Q�"� C�5QN�.�]b�J�'<��.ۣ�:̻�ϖ�q%�*(���f�7��� 3��n���HV�u}�3�h�ђ}貱�mb���Z��d�o�Zū��o�F98��$��(����j\
��<�7qڞ�5�������n'y7h��59=�Ə0��ė�+���M�!�S���'��n�C�J���C#״����09��@��J�}g4��� 4�\��O@={>�RrS+8�b!��F�i�3Q���ZbH�?}�3�$�}� @ pb�\�j�:�n�b�-�Y%�2�#z���վ���3��tBN��&Շ�K�̚=�<R���ޠ�w
��P7_�P�#Se`��B��z���i��j����x���(h�,L֜Bb�*������/���,.�8�_��U�=Q5owMӦ���V�0��0)e�xn�)o�;LZz�@�)��S�uNݫ^��L�A�O{z^�	])�W�`:�u��4>�YK�[0���sS���jk�ګ�PS�̓XuT�e�f5Ou+��p�ښ"g۵hUez8X�׃��6�6+�&�ǹA�c%�;V���3lbB�:��q[�cg��M����V��?���-ׁ�4V^�MZ�		��{��+���V��BDlb���;�L*�33��L�Y �f.NH4� R˝o���{��Kyb ��©q�V��Rc鑱�ٸ�H���d�0Şī�c>�a8�i�\�p�@����S���g6�I�A?���1� �>��@����֝R]����S��T�c�û?ʒ*kzX��Qa�Haj��\�`����6��Wޯ�'siM/���?�I��D�\D�{)���w�!7rR��]v<q`]�+�*x`X��Q�6��`P�����O`�EF:���=�#��[�(c��	�[�i��V�>d�'$$E�zڵc�ͅ9�:��7��^GfR�>���ԮX�c1�Op
*������<� !���������r��f��"�'�ds8��s�A
��z'3�3+71>*��.�/|�gt�uЌ�z�k*JǤ�OYf8�+P<=��`�OQ���F�5��J�p4ύ,�C���.�I5	e7x=����p�C05C�]��s �/3@<���D�Tr��}{ -�R ���,Yn���N���ԄϪ���<w�+Z����-�P����/on�[���_3z�ŏR�/���Q�A�,�G��A�wR���n�-��?ݐ���I��I�W�S�B���~A���3��fzŉLA�JT% m#�J�'��C%m"B�F�F�3޹"R���P.�/c�G�4>b{�����vo�ȝ�;�61F���3=�;8�,Dd��me����7�~�GY���4-k��U���d�QI��w�A�d��4/&p-0��3���-�0��½�v���Ȕ�^?THV�s�)���'�WM-^��~�K�bo֍����y&ԲSSGGE���G�^�aW�}+ � +�q��t���<'��E~�|KKA���)sB���+[�(����i�"	�m�!oU�^siW�bs�M�	��cg�~� �"���h8/�"2�ys'Z�4����NwC��E

J���mC�FW�b��n�����r��]
84�������3�i����\qip���%?�_6�G̀�y�EƱ�;�CvjSu_��/�e
\���Sq�,E�rkf��=N��)E���#[�^�9N�T�Lq�~e���L���Y�A��+�8��Ʒ?�I�+)7<T�����j����ʿ�H�av=I������U0�R&���]I߀�����8Ju="�/S�ł������n����nx�R�g���p�ֆ\��n=9gL����z��|[}��E��2�T:�u�z�D�*/�.�$���d?��$�C7�8eM˸0���@Zy��:�G�l'P�m�FtQ���̡�,�36&v�x���m��p���s�dX�-xN��D������/3����B|�Ȗ9HtLe�]B�{�T�)�x
x�
���d`5)��칍6�G��J]��Y�W����*���Z�@�������u�n<�~�&^���[�^�׆Mc�ش�J�����w��*�6�b����^Z����S78���t֨��f�7���/cR��� AД,h��c�E����ߴ2��������DD"�_�G����E��>F���%߹�_	E��nE�~q�+��^6�܌�]����L�#���xH�����:�H�+]$R!d�����j�ѨB&�iʽ������c.�S�����<���3+5��77��� �)I�m�4�ڱ�T����Xy�R&�	6����R��1WGW8�����b�і'���A>��ZVh`�1�T���=�r�%��m�t��֯���Md����O�;>OW�=�;�=!~ ��'��.薥�K����,0���;��3h>��f���y���� i�H!���H��E��o�ʁ҃`T��;e�ߦ��Rtm�v��EJ]��k7@?G�6>�X�s�~����`�����[�T����UK���//X�QI�)u|�^��iSa�:<6��$c�Ch�YG�+·BC;8�3X�0[�fa��:U5~!�9ʘ��i֡w'��0��pk����;!�?A{$]���=����
��
��9���M0�-����cc��ϟ"p���F�|F�ʆ2ׂ�z��<�_�Ύ��!�K:�X�Tр�B��-���6pCU�3��Ȅ*�����U��!��F_�t�=0U�뮬�*Q�t����i^��J�MTv�o5�e�B�(�s	�Wڶ�:Ii�S��"���Zf�t��� gc`����pH'b�������.ŰO��9CH5��F�CV�.leCٝ!pj�n�9I�ܦ{��@�D�%�_��]�V݈-�� �[�
I�Q����vsr��ӧN�Jl�m	�(�Q�	��'�^>q}��s=�%~��=�η���؀��><�����_e��e W�?�����)�q��2
�T�a
���+��?�`��6�C�p?�Ѓ����2͝�Pf݊6W��*���斳!U͸�&/�^��觵$�G�@g1c��/3�0�ou�g/&dIh;2���D�$�9�誹�[ԭ�N���x#i�x�:yB��r��g\Y�yq�� a�,��������N-Z�W�!O|*%k(&��#>�4<ң�,*D�u�=�;D\0󌫋퓟|J.PJTx��s�־������X�<Kf�EC������vۛ��C`���~��mV����zX�}-R��C)}7��w!Ro���X{6;�MW�c+2�Z�sR����.p����p��$�d�p�t)�B�E�UKv jF\i�\��d���XN�O�B�e�x�+��
$���ZL�	K���Q�������� �G��ك6��v%�D�$�쌱�G uQ�j���CX�f �;<b��"t]X�j0��A�;G�3��U�-w|�����cRŇ�*�k���tgG{�����u��17�\ՇBmT�5ti0�s��ಂ�#qi>c�T���Y����e�����.$�~��`u=0�h�7�d���Хl��;��'yX�Gs�CB%ȷ�k�sP�,;b���sv���4��A7��Ő�� rKOm��
�\�X*%���sO�Q^# /8ͤFo�H�!�9~�R�*j;��%X�ֆ�W7-��pRX���.����R�(���΢:g1q��L��� 	Q�~�-�=X��Fb��2�R��Hؙ�8��j�8���>��`Y�}"x�9��jr������s�M�%�B�y��	��.���_S��c,Q	OɑYv��f}wπ�4���@W�g���Z�Be"2n٢�fnj��[%�ﰦSK0��@TE�b���$<+���4��rbA�R���k���E�������F� Z���cU�[�rp-`�C��&h.x� �ӓ�}��#H��a��ND�Y�M���}M,d���L/Dt!� j_��F*�MU��9#�m&T��i
�I���G�1�@V���p��e�+��#��2�'Z������c$���U�FY;h�z)5��@
�������n�/�;��_�W{�@��>9�wOH���S� �����GߒN�h����2� ��z2XdM��f�
`�|�|��n�*�\�X0�4?��b�}H�pb0�Q��j���zXS6�H����#U1B�lw=q`a=΀o`)��/����>�`�32�����Z��A���%��帤�&Y�9D����ڇ�;V�0z���&�X}ws�t��-a�Lf���0C[t����!���,��:V<����y�=`���O��	������%�؋�1o#QR�ǂk�QUDbMa���ޗJ0Hq��e8B����5��A�~ҏ0����:�gj�>�3���r2���2	�	�XB���>4]�xr|g��N����T/ ����Ib�>��Y�^s͝ڰYC7),�:�\l{�Ǎd��n�vO�~�M7�U�	=���0�3Fw�sY2�ph�* o=ޥr����;�/�v."�����Q����<G.�D���1|[1�X���ts%�u�h,0�6����@�������;���z��H
o�6�(/��S�����|@nA����d@��p5:�^�4K�jw �����`�s1��4XS4]���ba��1[��ױ�X����,�j�-��)��B�@��A�0 /ڂ��%��t{�@{%���"�ų0�c�Q����G[Iy3������^mq�:VO�L�I?8�k��_�����a։������+�6������]��4���ƍ���
ʋh������T��n��4滛��	O��"�~+Y)6)Y4���F �O�g�.𳫽��9��def������2EN��;j�C P� �
��}/9}^�!� N0� �B���1:Dg�|<��z���
�Z۾OW� ����e^2�K�i4�3��g
*�e2 ��ܿɅ�/����B+���7f2G�R|tՌ��C֠5���-�ۆ�/�ob�?���Y�&5�PE[��;���iζ��:�D6��o�SO����c��f)9u��K��jϠq������x��Ў-��Z�X7n�Yr��zn�Q��%��\��">�������:GЈ��I��
�ͻ'j]���^Y`
����K2|�E��Z��W�����y�>�����l����)�f;ۯ~��]Y�osr��R�f��"o�OV����BD�
�+%���RA6QC�����#���&2�Smc�{d\�>m�̙�0R��L��0:��&L��t1��Ʀ}���s��@����2�*D<�3�g�H��М��-��Ť�����! �z��~ӵ}�K���8<2Nj�N�!㕞���Lp���,��@!���u����w�	�t��	�*:�(�g��p�X�!>�t���v�=���r*����j�V�r���,�ƅ��j��9%tu����-IY�O�\n�:����֘ >��ڙ]�ǞϠO��F�k<f8[/�a8sBJt4�����u�98'{ )�츌�:\��,��W��Y*���On�iC;���/']���W]���/�A�Sc�r=�� i�3��qҧ$��c"���x�$���������kԵo���Û�����JN��zE�iF�����߉v,�N�Yk�9A;�ֱ��00�Y�uV��m���ѣ���(��1�!�4�.��E��n��ӛ����+����	���)Aw_��K��ާ��	����wo���[��e�TE�7����:F�������*��2�M~T��<��~+�
x���7>�AQl�n+!G�Ҙ͔�x�n��C��Z�����ӛgF��[\ry�A��=um��k\�w,�]�2���%�'�\[:,Lu(2f�𔽧�7����+֕�۠0�b��m��}�mr� ���?D�1:\X	 mr*������o2J�`�ǹ&+��,qYNx<�c�Ҕ�����WI�������f�<ho��F=;Ǒ�s�͇2�$��!�Ϡ+����ѠQ��fߝqx���k~��BD��s�0>3��dh�>�&�>X�ކ�����u�^0<R3|��k�>��� �*j���]��1�~�i}�c��߃�Mg54'U8���u0eY�J�ng�;@L4H�&zT��/����#� �;k�X�	��Ԯ=l�m/iw�>=T�H0�'�8�{�[�{�	�p���=�e]R�l{܊�?+o�����������w_	ms�(�"��ƭ�{h5��Ħ�9��Z���N���/�����N�M��-�_�4"��b�k����wc�9�dvI�g�
��G�ۉ��+MI�Wg�jA[��I�4���*�7d{kF~����ϒ�$M@t�a;Q�w��.�����c��ӏ�`o�����/|}����Y�ÁP>�霵0�9��V�7��ᅣ�'���- ��� f삀}x�n����|>�u���
�g�X����%,z��6p)! d��6P�������p8x�?���-J|>�t0pi�oc�{)A=��oٞ3I�ӷX�
z���n�����bxfJ���U�G]��������G	2��C!|��]��%����a)R�g�T�g��� ��8Rq��wMv���Ӑ0���#|J�d�������G0�bq�J���j�U�ҵ��y�S��l����S�p�n��� k�Mg�^[RR��7����7<i���:/"ɊZ�r�AN؅M�]ψ�����?s�@��y��z�ڋC����Q�ҫ���tԓ�{�c�%�đ9�l*�߁%�7��� �kt�Ǭ9i��U`W�����k��9IUJ�
;Q��w?�t���A�0�:l'J><x��EY�{��x=c<U�D�E��8!h_���{�����P}�Z�R>_�����D����h����:�N�B>}�����	��h	�m��"T�Y�&d_�r	���o�>��Jŕ�#ܹS��B�����F}~�b����x����u��;��`��7���T��z�{^"4)w��9��f�M� ͧ���Ϧ��k�H(�C��3A'�?�� ��c�TW�]L�C��]q��m�U@��T*����	�C*�h��&�����e���i�k�ewr��p��!�#���x��sq��O�#�1�Mn����I�5���O�;�\_EM�YФN��{�W�A@���/T���0�C_1��^C`��L�Q�*�C�"7�[㵥(Rꢈ�.گ�K���h7�+e���g�Mܥ;rBw�i�!Fe���0�v�O:����N���nGBEٵ��=m�8�A��u�2�7]�h���Ps�H��ۏ^%}ͪw6f+z�����z|/�~��i��I/����tU�B&)������&uu��z����I!��N��C�zB���.��l�"����A����&R>�Zs���4N�ɡ���؞>O�����ݒλm6 �HѝxV#^]�����D�Q���,�%;�ǝ@�7WZ�e���w��}�[�j*`0Wy��}96,�º��C$�Gqۻ��n�E�.�I���[J���bsf~�wiz^�{�gx]��wt4�iN���?E%S-~�Q[sx�qX�S��͌.B��֕������.G�&P�ø���d�,H�`a��6�ʾe(��Kȇ+��l�0�M��y���h)��^��fǜ���ئ[7�$NߥQX����Uc�i˭��=�b�0+��@	k���� j����r���߅��kZƕ��;FS�\���ve:Z�K���0\F6�؄b����gҿ�n僶0CK6�o�����.rUE�=v$�_u�$�~��&�4|�,!+����	a���k���'�6�b�^�P��V�����T'I���Oљ �|S�9�"4lt�R�0���G@�m>ut�Ϛ��̌�@�Jr	�ģ�̌����vQ�+��@���J�`|��������ņ&��b6	�Ngvjx��o�]���5����
�Ud�/f3��>�����n�L��~�Q�����0�� �ߝX���m��vD��H�i.�?u�4_!r��1Ų���dv��I���/}��&>e�&�x�_�OE�Kz����;ii��&�f�q~�b�M�{�%��rӱ�B� G"����W��Z��DnV9jXEŝ�9��q�k��P��*��D�`��\�����|^�1'�͚�hx�[Pu½c"~t(����љ(R%Z� L|"�D������i$�g�T٬����Y�_Ld
�}����]j�DL�d�(>�M�}�����(�R�E����s�%���tmh�g)b��&s�����n��^@�I�o,_��L�n��x����HZ1n����և��␘7���f<J�7�Q�������OOOa��`e���t�v>^�D���==��������8"�c�Xȡ���rC�q��������gM���l�{��J�!M#�2�O���aJwܘ��<�o����nO��1���/%7���u`�fl(����}
@X�O�zh�&�-~&;�����D�����)n �V��:���Jز?�ظ��8���(Z򦣆͝���ڽ��Ĳf;{1�$�^s�مܯ[[s5��<-Jެ���v�BR\��-��\���Ѐ
�lCP���������H?�[(ɬ���ɔ���s�m�Vqs�u�3俭�^�"=�_��	�SupL���V���B�,5lD��\��OE)0u�H���i�T�f���C�@N����N�U"�j@,���e$�9���ܣ![�D��O,�g83�OK�Q�ks�ae�P���SS��;��߬yQ։�*�����w�iw4 ��{��f�e�7�K�	��̸���篮\�?^�{z6�M��I���n�#B�}>�h�]� 6��s��5�r�J,�f�#���1� ��K*�)V��(?/��������S�!�/m]s��9\BF5tr5=�#J��KXt�1Oܨ��RK���ye}�%�����jC�[t�xu!S�B�O���G�^���%��1&k���"����w��1��7 h�8~t�����w�s�/1�p#��z��M_CS������x-�t'����`�tT0�]�e��]-2��M�F9��~�cR�G��K����w��k��W����h�AV,��x1�����C``2�y6�,�F���ԋs3N�=.�Y����Qjl�	<���h�T� 5ۥQF^�����0E�V]ޜ�!���*_�������L�r����������h��BՌ�\�5���jk�+WV�"�#r'1B�(���j��G���-7#��4�i%�;�WP� ����B���ziZC/F�����l�+����Z#���5m��E��\�W%a:X�-H���ӧǲஸ�/Q褫݉��e(蘓�ѺE�3�꡷T�E�Ɂ�=��S���?��d�����g���{Pp|�>ɒ4z��3.쥰T@(�I��5�g�A�\g����2Yx�т����L���9-d,��M�]�,S]J��w���`̀A%֟��H���YJ���#�D�P�q�e�:icc>9S��c�'��c��p3�rIX ��~�?f�S����!�H��|��yր�A�=��B�>I���`��4���J/32�D	��m�`�R�c#g�����2��eͪ��4�����hI��߻������4�B/���K�-��9bcھ���M,$z��\$@�!O�5����a� U���Hbjqι��!�4;�.G�����&$0���b�$���΢���߷�U3�DTyx:"�`�Ǥ�W@x��l�D2�	�'av�	���ߡ�x�V�3G��C������4ԕ���)R��S�Fk��mj��Xo���5��8�~:Q��w_�T��cIY-,���}e�
���o���EX�)~�';�ԩjT�m�E����%�-T��Y
������<�:Q^6�� &��I�蔆��\�b��o *�x�#����r~�V��<M+RlɊ�nrE���]�N�ϙ�;W\G������hM?Ά*����R�GƊS`6�..p���×f t!Eյ�j�P��s�������MWB��@�������o��<�RHB�E�yJ���K��b�S�?��Խ���W�e^����o���<���w�M�;I %��o�$�E[���)}
3�o�k����Y�˙���2��z�W7��&�'�(���,Y�d��[^{l�Ml��ZS(��/
%��^�s��Z��Y��t���\�m^2?/j�;_��!	сg��]_cq�u�v9���9��/�_����<w��KĤU�����%	'��Q7/��v��.�l�����r$�
O,ƿ�>�a���N5�����;��`�2�BXn�E���/�`H�#y~��l[=��g��w�+�R��m��s���ߐ^��mxM����2�6��)1�]\�In�ِ�V�6Q��CU�ER%c�PDI�B�3�ȯ���AJ����ƴ�c�1��n4Y�AN��V���+5��Pg�͆Ӕ�1[Չ��\tL*K��X7'rFU��J53^r�9 B]XLn��:���[�����;�+�F��{�i+��|����m֟e>ɀ���FT��a_�z�n�:q6}��DE�%>���^�����oqn��7u�聗�2�\݆��-ٟ���7ᶾ��t�X���g3;����_��b�N�Q�=39P���Ȟ�F0�b��wS��:�b��4`p��1�IO3vn��l�n����v�a_b��Nf�k"��#o�F㿲d�*�M���W��Q�ԏdp�Y3�%��l��PQ����U1�7������(y^�X�	'��dqZ���*��:}e"N��Ai��������ib{o'��ԐsǍVe�3��4�2K4Q��t�����&4��K1�J2+����yJ
��b����������\E�%�?kc����=�1�J���b��q��1���$<%;��:� %�(�t�� N#�*O�7�>:�A��Ltq��k���|OJ�%"ƾ�F*K[Rd��.��'Gq��fXi��Ѝ����ؚB�&۹¤����J�$W��R����Z 1�<Y:����8�q�1��۬O?B���=�C?+��J�I�ꗹq�45�+�,�����׼2||�%S[*�꿡�L1�6Go�ξ�=I�gZ���~��o! )���:�{��o�%����Hy�����V���NZ?I��$!c!M�3�����9�m�J��}HB�H�ӄ����p���GmEb}0l�dK������ G]ŗA��"��(H�3| ����Or�$�c�o�}�׋wpa�9m%h�a���+�e����[���%��3�lfK��?�	*�m�HB{h:��J��b�����U�R����N�[吝໹�� �ʠ�5v�5���r���B��Lkes�_&�67�H|#���]���{�d����ޫ�Q�s� ��+y�Ʋ۹���5.��Oj�������v%��,�3C����S;M)mj�D�
n��-��1"2��cQ�rf�4(�(:�IՊ��H�Ț�D# �������~T��bDro�j��Zi�7.�_$fW�O�����U8Ӷ9��ޔ���x�C��*��蕸�`+髡�.�C��R@Z6U#��#F?��fK�Ѿb]����K���0�%}U�-'�u���Ԁ�l�L�ŎF}+��Ê��Rl�Iby��}ʎ�mðUŝ��ۈk5y݈�uulM�M97bOW�_2j�_/�8kDp�!P����M�Ǯ�Ӑ#/{�4F"f�m�WwkP05sa*������!Q�*�B�B���!�tUi����?t;p��N�N��c���֏Y��ƕkȩ�K�x8qcn�r3:\d!u	g��7�3 �����Rz!������b<Q�����.y1/�_�+Q�M��(<L b'�Q�����Ӿ��A�R���u�Nh���+o��.�HZј�����6�'|�ݷ=�.����>}��4Rѹ�lZ'���K@�P|�*��d\4e���|l�����D�8e�"�Fp���Z>^�x�(����Z�}���}�D�w�Pvv�m��e�86 �������[�L�J���E�<$����Q�	�?�iA8�c �t������Q���c���B*
���,Gw�S�R�����ڨ�|��+^�N���\�}�u_z��7Ǭ2X��K�DE�d:�5nW٤��7vZͪ.�����*9*^��R��f���n�G��L��r��hT�>p ^�*���37Ց;@�Ta�:���~�/�RF�����Y�#�iS ��e��̝
�DF���k/�~�?���$PA.����4ݎE܈�`N�ԭ�u���"��;A�7'�ϗ�0#����8a�T��u�"O��t�(�V��>[�*�]����{όh �*f�� �=�c���ld�MzR'�j�?W	�$NQ%�`�j#'G��S~\Z߰�F��|����˷ޞx;dIb�GG��$����"�|daT�3b�����VpC1�!mO:JK~��ӛU���jvd�'�u���$mcMj�_�PF]!�O�z�P��.˻K��-��Ц�8f�;�k����zD�I/��N���ͻP���X5�Pg�O���܁���^vJg4���*�'��Q
v����WN"L�Jڤ{��:������+g��of��I��R�v���O��Nm$�g����s=֟F�.��cQ�~�< ��,%(׋����q��6b����譝u�"��6ʈ�4��Ϣ���%%����Pq*�Ch�Qu�V���[�V���Ӂ!m�i�PI����'7�aYM����
�P����r��K�$8�ع��'����n)��~B�Y��T%�p�P1�����Xiv�Pt.��d�����ܱ�4��c��H=���׮�$V�/�kQ��=m���

�zN��>I`i��&��\uFj�wY�`�B�/dsG��xB����b��d��4�}ᵚw����Q���UR��D�c��x�*�g�ǩ��lRP��N�1�p�����=)`�=p�~�:��
�6�Tm�̜���q8o;��	��N�vסg��]r����~�%w?�r&�<�L�����v���-��]�����q�?���Y�8+Mx�8���*��A��ӻt�W9Ѽ�o?X���u0k�`P�v=�� c��I�V���.��h>n��й���<5��iկ>����x�!��%!�qR$��zr�ʈۤ�$>12���>T�-}MAc�7UW���V��KX���nR��Noܙ�O:�FU]�Y�T7>��0�c�ɼ,�D���&^�\�=��t�S���/���t�	!��Z��#�Q��ũ�u֣o�Z2�=�qyF-*K&�q�5���� �D1~ '&.l�=A��k�Dp��&��;&P��n��*��$�=]-�� ���������Ws�>�Q�a��؉���p�Ч˂+�ڛ��x��l��r�Ӑ���� ,;`�wbswvq^]k2��l�3�#^�3u:�t,6�#�3y�8���m�H���P"JD����[ZF(:��x�_�|tml���ֳ��l��t"�8�r�J4�A�1��4��I��g^/xntiJ��[|c��q�����b=���l1s���:)��}\�S��	C���E�y�܀�8^5d��M�h<�Ο�^T���-	��������n��/��7}�S�_�OT|�M�P��kWq��Qp:�LR&D�3 �C*b�Z���Z�pe������I�	d&�o��N)�M��嵼"5�G�Ǎ�"o_�-��_���E�v�q-ɀ5�IVjh�5�؂��:�&��a������[�J>6�ɠ����/{�eS~p��c~��<p�4�f��wT����v��Mq6snt���Đ]\_�\�t���L�^� o
K�����.\D��u�f!ĕ��	f>|y�����C�هmK��FF��\�@��n~C�{�V�k���y��q)y����8�v��'&.G���:�-u�.���Wڐp�~��1���Ǿj�>4���DeX�ؚ�O�/����7 �d2�C�ʯpA�x2רS{��%��B��N�A��|s4��S.&r�n���/(;$�ŶF; H���.ڄ��Q�5b�>��PRΚm_P�d�-`�g����X�'�н`���:��/�0U��i��E���0�K��h���� (Q����W��7�W�tI���*�up��<��4����a:�UI<8"�)?M���1$��`Y8��t�0z��#�D�*s�9j���sb��Z�Vi+�E� �<�?�"&2��s�yÚ��̴1����cq�2B<�,��v'ɿ]��cz��{L����S$
Զ3z�j'ń.��y�Z�؟_��ZJ9��?��H���Κ��/���$���&-��D\�Ih]P?>fk�sv�n�.����O�KGa!f�|P�����ͧ@:�y��Yq&�SFu�⶟����<����Z�%�))$)�G`r���R5��&=����T��P% 'P���$D7��������s^������*R��b��t,G.`ĉ~��ն��{Yy���~�=��P����Qԋ��G hDf��z鹥���V�8灓��;/�t��n����A'�Z^�"��-VnP��\�x���A��%���p6����ʆ�N,�'�ɜʔ�9�@��4?�0 �����}(G��M�Q����m������Xjnn!����g�v�'��{��-+9U���U��Ụ$�G��M�k�"FU�B��ԝ��X�ʀ(�&�twIw�4K�t/)�(�*�t��%��)H.!�!�]�����}���Μ9s���sͭ��vDM@Y9��*&�ޑ'�cXCoax�/m����<�+�21i�ɸ:î����5{*=�ٱTd��p:��p雃� �l���LLբt����"h��l1��x�8m���>�j��d��e�^��B�`Z77O�Y�P����q��%w� �Wa��co@�0ĳ]m����Q�\��v��R8޿ճ \���4a���ꏢ��x��fC���oW?��
�T��K-�V^d*��$yfF;���E�+�xا.4J�Jj;���E���y,�ky3������а��X�P1)���$�+)�-��5Q�G���=E�_HgS7���ī[I�OB�����;7�|]ͽz�?z��R�Y�o���O�S���/�����vy�xX��E�h(�>�/�ˬ��Y3�z��K�ZWn�ra6C�b?�+G�h�q��m:�~ 3���ʵ1���=�Y�_�����]<Ҝ���j-y��/�?R��X*����ɻ�1��|����dK�m�>0>o�k��ٳd��l�s%�������eM�/���X��&]����a��"Ҽ��1|k�."�_� �ڦ���8���!&ڰ,lYy�����N�>��1�2����-��	=QF&��C�dޮ�S�ݪ���Fh�q1��ŋ[q���"�ŏ�`a~��6��_WrD4,x�D�A��6�#��[��"�F�M���������X����Fb��e5C�ܝ��}���}�7h��H��J̦�T~��=ɗU�=��D�]�'��:�@ҟy
����w���f��ah���RS��{Jm��@Oz�Mh�;�*i��M���43;��]s�����`��K�����QU/��O�!]6c�����s�HyO���()x�FϢ^�������I���Y����W@��q���`�%��eQ�pOYe���=06��-8OibX�{�cs�ֽ3U�'�Z�<�k�M]H�ؙ�~�3����+��3��XǠ,�z�Y��oX�N�V+�G�ɏ��]?w���\�W�g(V��?���bR��-�jq_S�ψE�_sP���qgz����O-+V�و��"j�����j6�36#��oC���ɍg��TC�)����9�2����o�%9)�"n��@�)�Jm�h�GKV`��؆����$C_�~*`*R�2Pr�q)P$�������t)/Ui<M�D��Ttk�������1�%g�������m�&�k�Ɵ���5�8a���z�	r�9��9��q>���_��G�O�Yl�TT{-*�䃘wsFFJA�s��0>��L�K?S���B�
��K������n���s�:�R���r��O��g��, �Ijc���0�����Y������\.��
C��k���K&��R�s�znͧ&[����S@�F��#ȴ���xվ���n��5�D�z�G&/)�kX�s8&�=���/*M=�@C(۫rځ��bN}�ykƅ�d�Ikf�Пy�L�]B��`m�'���j97� �Z9q��7��Ԓ	K�x���D}�>�����wм�Ϙ�t8�����=�u�B倮�o"�g(��wCP#���Y|�F���@��0�XK�BA�cLgl�v��#kJ�$��։o�>�[��#��,�B(�y�I��>Kz���3�С�,���̂z�|���kkW1�#N�]ѩ�{�t�)�>���:}�R���8����G� $�J��<��'���H�0uˌ�����48��?�]j���.c ������K����O�_���:3�tz?�j�NA�'H��j��� ������!g�qXc�Ά��	�1���9���F�PU��������I׮V�Mx����F�����)1��A�I�գJ<�T�P\(�9X:+6����7�faD#�������0�ȇ�	j}^�6�[_���]��FƏӷ��&ԝn����Y)Y����?ڙ"4��mB���}6��0h)�	Q;ߎG�d%"��#�?�Ty���� D���H�'���1Qr�L���
�Y���2�i�0��Ev���T����Jo�b����<]�����:xFL�oB�<nm�B��vl������3��<���'`|H �S�_���[��I=tA���V��n�����)��$�E2)���a��}HpT��q1Z�N.H�ܺd�ehWBŤG<r�	WYS�I��2������K��{�P�b�H�Ӂ��dI�s�"���'^��_�<������L�(SI��F��12�����\3^����+��b�?E�x j�S��Ӥ������8\�,کJu�z%������L㪅�U����+o������2X��Y7c�kv��/RN�����#C?p�Z���eF�oa��.,]���&7H�PB�Ȭc��^��F�pS� ���P#�gdw9h]�l&1~F4u_�kNї8HT�2{��Ah�>�,�[G�Y~;r�H��A�66F(��uM�I���%�����$B�+7.�:�פ�3�$��a��
Ϸy)Y=\��:m]Xz�#���#� ����s�\ܙㅁ��ʙ?z��s��-�\��Ek<9��Z�y�w���������y�s{uY�����UJe�𲹇m4�c�QN==�w2�yr�"�?�No��8�s�.��`������	E6�">�(�.���l�P���&�֓��^C�m�&-�n�	��X��4�M��NbH���yh�,~f��nxtz�]D�`e�-֒�im���v�aʶ���\��~h����╃�<�X�T~���;R��hv�KI��zI�J�!Je�4֘׍�@dg��Q�B�?w �'�A��}8׫mğ"��e�mА�8�sѦ(�0@��s��~��P}L�3cЀި�+)��oV-x��D��	���������cG�S1Y�[E�Tx_��[ᓫ4�/�*`�2d��I���\c�J��� �����d da%Qj�R��w_o�tR?�rDv��Y �R~��!���ʆF���7�y3��є~h���Y� �O����t��K�$tK PZ򗝩�)$b�������<�T!��\��t����El�w�?�{������!2���Ԇ����tQ���_��c�iיHr~��W�#3엘�O*���Z��9źUo������PeHW�?x�{�g4Qo� H�|m~0@/BsP?�fooO�B��� D�1"i|��m��нH|�!T�G;Ɖ]��o�6^q
���>!���3r����Rֈ7Q�O��ت��0�Q����_�J~�{�~뾙ԇ��￨I:gp.����a��q��&n����g������|���UpP�[�8�DN{$47V�/���bָE9~�1R��p��q���K���0L'���x�t�)-��W�W���ſ涗���ώK�v�S<�5iE���7��c$�����f/�5W�Tx;P���7Ԁ�'��E��(x9[ �	������dq{E�ׁ�+�B�N����<^?�Z����֢������J�V-�g�|����Q�F�/�$�-�/�v3`X(˟ZT*��|2�F��u��� N�)A�U����rU�1q��
6���M�N��
E.��'��t��bBe�4C��z�^'�6h�Rk�HZ�:�/$U�z���=�tH���j��@8@�5D��/���+��� �G��Ĕ����i�����Q�13�mfz�l�UV)խ7�h�&&et5MH�i�R�T�z^��,��|C���In Z��o�E��^���0��P+��d��7Z*��cI�i�0���:��+[{?\̯�m���^B�h�W�s��4G����Ph���:O���zuYu{���oq��Vu������О��f±(�hn�q�����A�����*���p����'^�]����R?`5	����6i�T�*k�aY�4�
xj��y�B�N	�w}>��Z`iT}C����Ր��wxPv�E�q�3��b��P�<��k���("4UU�(��#LCt�~���4��$�{+q\��㜰��m����P��I���k���θy�vj�M����dT簀��F�ۇ0Muq"��l1dc�2:��+H�*���C�|��9Ŭ�g�,7���%����m ��)��g(Qv�1��J���A�X@�ڦi���{���?ˡ%��8b�K�i������Ikȫ=/��M=��4Ϯ^�B�)Y�qq��*��@�,�~�����q6��y[^�����E�˳Ex��&�*�z�kXh��S�d�UYK-��"a�o6g�
9�	J�:	^}`e�bh�=Mk���������V�2W<������:���*̘�'�`��@�eO�k����v�����,���y��A��E�����%n	nQ㥹�Z�4ir�o�ڰ�6��ل��n��?I;�n�X �������]a^� �%�X4�Dά�L,i�X��1�4����gE����'�~���==&����&���ѐ��tG>���V-ףm2\ �ú��t�HB'����
l�/����,��'����T�'iH#>_�?���o�p�]ЮK?~�p;�S1&�#���U[���t��Y��퉳q�� ����F�Kh���g� ��M������3i��h|q���l�4�zm�w3Áv�=�4��,D�������K�z������	�(����?Pp����k��HM�^��]���EͩK6*88,9r^2��J��]�y9�o��jΊ��0Q;�����y`���G�QK^���8���}����,�x��wG�
�z;���!Mv���ǿ~n�ҙdY���qU�Љ���N�G],�L���DI[kP�&����yg���6��mwX�0v ��]_X4�'�ď<)�p������W:9%<�'�d�5�YhI�F�g�Q2���U-��"�k�I��ե�h��&kǞ��R[�J�Ͻnx��2�Ć�6(a	~L���~kǍ�J��כ�L���r���M[�H�y�" �5*�.uF��������`)���
���`KU��υ=[T���� �"s�С�Xb�|\�vX�~���5�޳���%j����p��4|�Ov>=���x!e �f���t���9�~�.����4C�\��#T�#4�~N�7w��Y�`82WfYVKG|LE��Ѥ��Ѵ#�W�IAĕf�(��mV����
K�y��_:bl:�x��e�|�B��,�8��o>9yEV.V����#;1����0�$����K�t�����~
 jN� `Fj�OShjD�{j~��#[���<��u܎XAa�p9�>os��=�(K� -�M�.j�L~�k$E�}�#�|���\�Z	�h�ᔐ���h8�����d�<��jך���=0E��4�c�J3��،��߆e��c�~NF����YH=м�i�Ҿ�2rҶQT{�і�2ׯ�Mx8ZjJh��d�	[�E� �&E�M'*��b�a������&I����(����H�^�نoh�4O���.�`(-D����F�W��aD2�lv�aZ�GK�Y;:2���?T��&�|����L�U��ʍم�œ��I�%��>�{��!��<F���Gp�����"~h���i������^��t��fu\���v���#�*\\�p���B�P;>*�.ӍTf��>.��]�p��){Ԫ�X����un�Wܝ���j��E���ऋ�&R�8�2:���%x��0D�I��yP�`[ɸ���H\�����Q@"l�܏�w�L
�2��Qfi˄6���_�\*6V6[�(P(j��}��m��Ȱ\bNA�H�������٭��	���pX CpQ�L�[�oN7��@�+�or�~�ܕW����\���U]I�L''5Bb����m`OU���4��H���
�~�\�O��'/0p���(c[�s[����/�h��9S?��J���.k��S:ʱs��Ʊcg���.w�M��7Ī�	9xC�(�M�zد�Y8��:��{��(?Y����*O�}�~=xc��6ֳ���j��N�9�=��a�����ԋ��F�~��q�<�:I��P�e�`5�}�t��>�LÉ�9ԣ6�ʰ����?��#�~,%)9w	ۡ���^pI�U;!\�Q��y4@�S	sH�i����O�U�����t\��MN���?��C�S�^���?5�ߝ��g�٧�/�C�
Z{�`@���T*�w�,E��9B`1�y^�����N�=^MH�,��m⩲��G��*�ө��ύ��0� b�1�̊Ruapf������D�ԗ(@�m8u;�Xf6`*���:W��b�y,���2d녝���mC=�l�bP��R�5r5Q�"AX��;�٨��>ʭ�Z��6ڠK��P&��m�܇�{�Ω]��r�^�0д��s�`&�j}2��Mg'�#l��1d>0�)8��
a�K�I�{���#$J�v<��'"��P`ٵ���Y�t�7S6�ŉ����[
��d�`�T�*�6ͳ��f@�|���:N9�Vo#�kS�w��[ʉ�^���Ȟ�&�Kg>�Et��?S�`���@uT�>�_�%��0�M�'�9*� �3-j�=�"�����)�V5�:�R�Uy��4h�~p2 ;�s�mW���� �S2���&�_�Đ���ٍ�r���R�C��o߬M_,��NǴ�tTif*T��"]�'��c�ʄ�y;I� X+V��j�McO)w�+?�?��/vE�-�Xrs��5���8#���{��2@�D6�T��p]b���kp3�N�[\]�|�>�j=Yt�n� y��­b%��ת��Y�$�Jf���Mo�wEH3�-��I ds�`c �g�!/�Uv,�H��Du{��~���?����v��� Т��C6���Q�G�e�f@��F���M)���a略}��?=�g����W�g&������nЉ�vӷ��ⶳ]��:!}� W�Q��+q=��#U �x�?��@#���B`����Dl��J�=M��Ê1�3��7��^*p��T�b���P;~~x��%7,�=�q��9�vÁM�K�U���/Y�<���]��Dh�rߏrh�H\�L�Ҁn�1 `�m�ܼN9 d�Wiu�	<+n�n�2��|�B��=@�ff	�6��đrէ�ɗ�JA�h������)�^ .���2�Q��H\�"�2k;{�ይ��X����C���L"��v�h@��|��Nɍ��eG��#�e���f~R/@�����jy8������
O�Av�&X(���ԄK��t��%���d�ܜQ�T��4(b��/tv��c@-��1QV��3��^>Q���ZBa ס���~�L���h���J����q{�c!�]�i�_0a�d�#%�>�^�.mcҨ��￫�3�~Mi��}.�r����hD����tڢ/�H�ӣ�g$��Ҟm�

�"�d�nq%��䓣5����$��I���&Y�y�r�n߾���ÓN!�5��@/ɷ������	C�8Y�)>��R���%�� �yN�uL_gj!��>%�9�D�D�Z����F�O��A)�n�B)-o�0�s��U^�ٟ��%~Og���b���9sU��7�u�VG�_��cc�L
��+q�{�}������x6?q�ڙ���MmsRz_��8G��>ڰ�ys{Q�=i����恓�iO���<�h��V'E�2�/���)��t��Q�̌���'�ט�J�����:��C�+��]`�g�!��\/��fjeEw�ǌ�m�*V;��)����t:!��m'��Vp�l���tv|��ɥ�B��]쮚a«��	�,�����xs�,��9�f�?���(��l��9!�Tl5�k�L!�U&���ɢAjg�K��fs�
W���A��OH��֙1�C����ڀ�rq���os��ɑq����t[_��B�~K\��g������
L"�Zrb��ïU�ߌe���L�D��~��k��GԀ�Ta�ђJ�@B {e���a���*A2刺�����9����d���'"���!Y�gsi�����t8 ��һ�1s^�<�ſʅȼ�᭩R�-��[Uba�J�~�*CF�P���ߌ
B����m<v����d�+DF��;+�p��u?�]������w.��s�j�����(`*�T�J��t�hU�`B|v����V;q�2w��>U�.���d�BN��"/OGL���>��m�eGm����bb�v~��ʤ�6L�|�zw���f��^E�Ʋ;�]Z~�1�2a�F1�v����}���:�[�_fu���x�i�uW��%{�	�H\q�o��tXv��2�C���P��PD��]-�������M��x4�m4�Qd/D���_w��ާ Cuk��5��|���,�`���)[�ђe��=#���{��`;/�n����H�����%�{x,�	L�)s��|͊�O�U]�0�M~�c[��w�ۦ���K��z?�]�L�a����+r��vio@���!i�2�`VR��_�/G�� K����PG�KJ�(M��� �R�V��08*��	�y:8�?_M��D��6W���MT�0�~��@%��-��Y��Lզn�@���̦��e�&@T�'ǣ9��-�7:��sj'I�u�t��f�����IPrS&��=~����!�8��G�R��{vΣV��qݭc���)@98$̬�X��w�ZP�a{�
K��Ki�H�r��հ��I�5=h���֮Tn�]Ѡ�t0�{�.�at˜:<�I�KGp��`���v#S��'?���������I��6i����+�['�"O��E[��$�D�X�zw�������1�Wġ-@�0f�xᦷ���G�4� N�(�A�aE�̯\�Js�.��iV��'�Z�	�)
V�?�M��y1FM���:m�w*�7�jh�yy!r"1�Q`)�N NQ�Iw�
�l�̯��Sj�r���0�����ј���yLr.f���`-V�@HO�}ϊK�o��R����7.��'�@YLE�%E��}�@�E?�V�� R&S�X/|X�ي6��Z��������f;3ʇ����Të��A|�|~���7��l;�z��Ks�8�0X�G�G�����=Wv�hJJ)��K��3���gV��i��ƛ{�<������u������X�D�wa�3x�k��εbsG+J.҅��[_@�gy�:�j]Nw_��_~L��UJjCR���]<(���ܣ�q�"B��3X �o�Қ=:eY[�H7� QK�(�M��צ
{��_;�=��iF�c�+u��je��!q
_i�F*z��J��+��C�u�e��;���H`���v����v�pk�N	����d�"8�;޽���h���P`�@�w뚀^=*�F( ��E�p������@6���giT���,���@�(�Pgފ��{������=�`��#��S�%"��|�$�O�ts�<����JYΒ���BN��<��ث�P�2���i:ھ�"e��QĈ	b����Bڟ�y�]=P���_�I)b���	�v����bBO&�tD>&�����LL���X��6�����@�_�R�y�[�D4���G��cg	�z��1���m~����jt���K�{i�0�����x=&�1�w4B$"#L�΍!��wgnZԥ�2�*Bq�s���,T����G�l}aW�1�w�����}(Y�4r}�k(��iV�9����3�a~���EMF��,P�]����^�z���4��(l{�ꇏ��}�'�p��B{�F^u��6���������2�<�%�/���W7�| �>Q�-�|XBb���o c�Q��.��Tg�DaZ�RY�1D-�^,c;Ƭ
ǜ�Yn�w����JU�G��������y�U5B�Io�6�q�������r�aj����s�),T?�~�щGS/\v�>E-BP�	�k|s6,���JZm[.&�7H3���F���v��G�q�_W�*�
���?��"�#)�|h�� �J7���,b0�M�Bw�UP�.]�i]0��ο~��D�Z��|�]����D(��)>P�G
��"��p��_cgяG��Mxa$n*����zx
��)�!=^�Iť�N�ps����;io�H/J� if�=�Iߧ�E6>��!@$�݊��*��M��K^����Ѯq�SÕ���W�eK�S"�{x��������*�^{O)���gv}s��7T����1/����Cu�s� 3�]qzUdO��^�ح_�����������W*�"����+o��[�Ia+��Z�sM/���U� R��b��_�N!2!B�^�y�0:�����4��lg�^8�،��I����L�)�տ"}J�Y!�?�i�Yؿ���#h�'	�I�\�7��(o�Gj��Q�m�%��pin�}J¯��bp����1�i��0�<�-�.s����J����lK�~5�B�8��e��Գ�#Ɩ?k>\q��l�ˁ��D,�( ��)�+CO	רf-R��oK�#~Aә���'^-�cNC#��_��"\�T])��#E�Ҡ${N���u&�)n��6��I ��t�\��8Mu�JP�a�y��2W�7@̇����}XB����k�z����3?_���9�"v%W$f>t�&�+��鳚�'��9w�L�`�m�kɸ%��PL_��,@��C $��0#��g���zai��XML���O�:I��tP�dЬ�Xk�0�yw��}5��5�u'�G?�z
.�{p�]��n�n�hl�$j����R��^��l�v�srd��'�\����O��.lε1�Ζ�w�{qo�4������	��������/��s�|1���9�黇6�Cg�:!���U�p0qL�e�a��<u��_v�j���C����x�-�ˮI�]�̎,$��f<{��w����W�������,c�a
������we��
�*��?�Kp���]m�� .u��V�X�s�N�e��k�6��[x�t����pSS�7,,�����l��Q���mwb��\�"��f�6��	�*�N��(c�7��,������Ph�Oz��@�䬛��%��#���_[}�̜�B�3
�ds�r�Ģ(S��L�\��C:Y2i�«�`z�!����)+7�-s�sy
v������7�2���M��T)XM���_��!��
��E�����<�P�����������#���	a��=����^�UG�����Z
��]��E[��ӝ�a����r���Iv#3��{��iy8Brח�le��&�*����dHO���������\^����[�IzDi|UE�<�o���u?b(���w7���!���ǖa�f?~��h�H���!�`�i����\��PC����g,�N��<��[�wD1�|�E6�U��,�Mu{]��s�,��~ؚ�P�KV�;�,)z�(�y�Gq��	�� �KM��6`�D��4`��I^b�4x����7����;��z�����b-z�p�j;UqIrYp/{.n
[����}xc��f{ pD�ޜ�͔���(�)1�r� ����[��W���ص;�*��c},�57�ݶr����D("_,	ZTo��#�1��g�A볼H�ď@�Q��GQ�A����1�e��?�E�8�#/�T9�\�x��CnkXd���-u܈-.Zx���U؅�^q��<���Q��v ��!�s*�hdK�1_@I�#�ВRa��>�җd0�F�;��F������c�-	�-�?�FA��R�x�jb��:F<xyP��@z�QG�r��kܷ����6��i�,x�:h@'��C�<qV1m��fU�h��yy�suȽ�t�k@l�|�	<Y�b�.��c�\;�m�۰�ˊ��b'��R��E�����v9��2��4l�a1 ���D��t�F��+nER�[�ȡ5�LT/qN���x_ǃ��B�f�NJ�{�Z��Y�����M�_�[��@��n{���(g{�pʦOt>��6��Sgs���U�6��G3���%,�e ���f���Ƃh�!��xק���d�kxma�<�!�ES��"?������r�7�t	E/f� ����{�'y��s�b)����뾵�Ja�}�/0�D	bG=��o�@* �|/�}�B�UX����_6"&�atsGl���:�� ����J�;�X�d�ZvF���(Tɫ��+_���B�w\6G8M���p�����u���>3�W�g�/��~�3���}*���@��o:���1�"�G"�q�j5����'i�Q�w�c�=�]�ߴ}�2���[c�o���'7��?4-���5O$�׉!��$&BjF��F�	�HFK���`�f;|!9�ؤ2�3=�_���gǉ��B�m{w��x�̆�$Sլ�9��r��1�-X�r��K)yb��j��s�[(qr?u^5�¾�x�u��Ĺ���XAP=�<����N-7~3������m�\�b�RZn�d$��5Q\��QJWMV�⧬͍��ֆv���JuQ�)��[����ݭvn�43i\צI��������<��.;
��b������j�5�����K�TD��1��q5F7� þ���Q�񀘃�s�����z��Z�fx����C�>O����a�y��������c�L��r����\$1�[jY�y�k�n$���Xǀ��)X��ꏰ#k�`�mmy~�}��m+�Qi+���.��x��WZn��'��欶��+㼂�3��K�G��'�>�`�p�������lW�<o�<�8���1�ʛ�<~6x�b�3s���(<�H{�M�z̄���.��y�����мG-�ϻ���wL%7���A�ӘO���%]�IW�U�ŧ�1�/	*BM�F,X.��!Y������H-J���ob�o��^]�S).�N��+P���p�A-�זǒI��P\������,������Y�+BP�Ԏ�v-��"W�L?����Q?�w���3�m�RXK�N������K=�xH(+�"D�Tx%I1������r�3�a����_���V9ѮީSh��"TR���p�@�8xS��׸�����9���!��ͯ��Цj�z�_]��%0sU(��̬ѕZ��+Ĕ0y<�*��h�w BoR��vI��]9�Q�8�
(uz���_
4���T�|��_ �5un��B�?-�ힱ�*KdP�\���L �����'dx,UP���>A�p�!�g;[��죝�q�NǕ8M��)�2����h�F'f�4��/�t�H TU*��4�����.k�;sC$ӛﵻ��(��zhX����_:��������G�L����U!�-���j'�.�$����_�D[$zҙ?���a�����>�7d�����h}́�w{3F�b>�(9�8����@f��wJ}���&[)�(%�8R/#�))&�?�\�;����*��ǳ����"z�"r���1{���J��SfE4J3��������տ��H�ˍ{���kE��m#�]�2DQ(�?�.�|���R�<����p����')�q����k��8w<��H����C��ई�+
i��	
��.�=�O(��R��x7&0W�����*����|���و��¼�S��u��'G+���zg|O����N�FI`cmaJ��/iR4v�	�5..T���/�G��������EQJ��͛>J\�S��0Ur9fc��,�ln=͕���HRG=h��M�8��� G�=Ad�$��*����QrO�H͖W��O������a�l Э�+�GM����
�� J2�b憓��1%�Y2�e*4���3H�����=���e�NBOu|h�$��<�4o���*�:P��k�����Ė�D! k�FV�S�7��D�_]�\^�L��j�M�P�+[�*_D�'#�`]�"��i@Ӂ9)��o ǟ��%�C�+4s5xtSu�9A|A� w�HK�<3�	=�,U�<pi��a�V��#z��}p ��s��E�XZD% +����u|p���֦��˧�4j�Z���a�hV�)�-�=�>�^5����.��-ԯ|�lm{8�C�z;�g����ӟ;���M\����P��|-X2.��O��&��#�f<�bz
`��������o�{���m7�����jP�?\fǶ�dYT��ضgR�dK��2~Z�g�&�����U_!��z��Bp�iMː��:[9K����뻹����vW�0<�N����}F���"���	�f�]��Ƣl�j�>Z���!̜u^��U�;\�ڕ	N{�T��M.
(�S����N�5����{y���O3[�_��@�V\�{Q�*�6hi��n��*~��L# ���jX�m���(��(_��*�-����hw�A��r|J._��?��� �I��ϔ��x	����y���g/=9+-�.�ҍP�U���7I��
���5���T�(�s�O��l��dQ.��ޘ(��(씡�o'�����t���"7�-���a%>|����GF̦'n������`Ï�iR^�>���R"�x��)|����E{���+��(��{��|�㴩��4�ꛙg����f{$9MM�������~���:"eD�R;+F�$5k�7jv�|2��B���+Gξt��eb�,�5����0
9�/E�Nƫ$b�n�7t�w{�5�D�+�ʭ(�҅�. ��>(]��O�>cy~4�s4.�(�\�F}3`����#  ���;ƶQ>i���܂_1R������ �8	�}7�!�gr���a���$��:z���Z5:cb�Ct��$��)����h�	���X���1?q�
�ǘ�����ݰ��H]b%Y�E�/"uZ�]���7j��F�1p=o	�FJa�J۝�/��)����D(�;wv��z�fO=e��(����m���^��~�eY�!q��׈VXvuVV0�,�/+&d�"+&�u4?[$lI��x��nxU�p�6��V��o�L�"��%2�]1�w�.8�=K=0-�P�L�zJ&6^��<^����M���ڿ+��*�u���C暶�"W+�5W�����F��<���$Wt��3�ǯ]�f>��ȦeP7�
�9�F��!]��ŋ�H���Л?�p�h�M7tb�@FN{�Y�,e��ؽ������û��!���5�Ǚ�S?ӏ���u1O-��/���Qg���!���$��=��)�(�ߠ�i��¨@C��f�~��ź{zW�)9�^m�\��Z,�;nz�V{����S�Ym��j�����l�o>��	�zαOvu/9�f��ihG��H���x��wS���	��#A�����\F����O�K6�)aM�Q�203Rk=�&��TG��o��n�s(�_��G
]<C�_��y�d�(ז������`��ضIƏUF��*̝Qy���"d��4h��;�w���2BB����?*E+�z��jN-E�(gڊ�� U�IL����D���4��P̼�������k~����9�ۯS��n��C��CS���+u�uG�T��%;CE��e��,fbb����������8`����q\��U���c�����x�o�}�'((�g��陣A�����dڝ�b�"M�ޗ�t���x�M�U�4]�
�a����y�qS�R��j}��#N�Lm�l��6���D�Į�9��1	��g��f�!���2�n|{ik�G�KݶVJ��*ɍgN��X?��L'���)�ٵ��aicP4�c��=�`���%�md�}y���e�q�����F���a�b4e ��>���zO�3�m���&��,�?�����0������>�p�X�חtn��0��o��W޽�>��۞�o���`��#kNGi%�L�5%+cun{Q�o���1GyŚ�3��g���Hɢ��#JU;{4Y�g�r��Ph+��͔�+7S2N����O�:`85�!R3�N���N_u���P@����c7���3��h�r�7`�V��VB���0�Fy
aL�oZ�2�]˟�y'eQl�)��ɣ��)hŅ
�#2&~i&.�~E���>��~�J}h��3�f���Ł^��N"޷I���RyPl�OC�x�����p}}�,�|3`j'=8�?�ֳ������ߙm��^��p����= �H�o6��}���z�h"+=���H�B9��NG��3�iU��peI|���*�	�|j��D�VҚpaO�T$ATJ�C�ʏ�u(�F�i���]�W�;o+8f)��ҼG)�	�B8��N�� N$�[��E�����sh���@��-|!z�tL���P)��Q+
�y�{� ��`�.�r�Ĩ<x�:��)u::����vM�X=��'��jӎ�����n��K�;�ރ���f���I-�Ѯ	 !��Ƽ�D>�LK.��y/��8�m���y�~��uI)�4*�&'C5��(�C�E�X��4g8Vd�	�fS�r�e���^�x�J�������~4��F�إ�dۂ��W�u���u�J�1b׌�j�ޡ���ڥA�U��Y;V�{���M�PEJ�U��m��֫��ཿ��=�9�9���s��Xs-2�$��0��ߝ�Y�OԬ���]4�2pU��sU��AB�����EzR�s�ȋ���L��9�G�)s7�0q��19��O��s���ޠ�S�����(��a؉i>��h)�˩�7,.a9��\܇9n
�򅦎��S��6G:���OL���2��쯇���m'�wDhK�fj�u,�k�����@uZcэ��͔�8�W!����3a�q��n�����.�����P�J	a�����z�]�)����#�i	A�Y˵��oLC��Z�6AE�	j]���J n��3v�=LK�謁Z��OV���V������}P7�Rtwn_X������_hi>{@�XBdNO��ߟ�!I��_S+bƞ¹�~���ֳ�9R$!��]l�-�����!,�E��BT�W�"\0uP���ƕÝ9�~Cܺ�V��#��T�g���~��EKJ�^�%TiK��AL���|�[�����y��Vk���.k_�;�&x���,s�x�̗f��ިj7+p~-�k%5xCݻJl��m�0���6�˦磓W�X	)b&2�l��ã
\a�]�Z2�K����i�M�����e����L�h��r| ��iT�Q���"f���%'��,c���F�^cH|�T��?�����`�zOnFْ�X���Gh�� �s#:��O��A|5a�G�N�dEj�l)���,/���;��=t��]��x57�57�ة���(_K���M�e�hGȋ���~��{'��Ϸ0�sױ���ݻ���;ޑ��-07��z>/�Lx�1�����i�	�&�-D��_����E��� ��Rty�����n�':�p��Z���u{��*��`_�(*�/�&uQ�͋�l$���Q�Dft�/��|�?�D-���%=�$�/�"i�����CF0&�ac��"����ê���:?ņ���3���VĄ�̀�u �r��^
���j�V��??���䪯U �/UM$h?r;��AR�ka醗;�5�-���A+K���r�4t��@Y����k��<&p0'�����E�金1����6m-�ap���r���ӷ[����_�<2{j���	�De6qN꺎��h�I���}���=� B��]$����o]E�hF���R_�i4����;��Rȥ��2�G�{�j��` �2�0��x�tJ�z� Z���h����H�����i�t娾�ߏW`�^U�v�K2>۔�Z6����V6���)������lZ��r�?Jˌ���I��򂩼d�9�fÁ/�t��sgȗ&��y���>�щ� �����]�,��|#���0���!\؅�@��A���v�"D��,>η���l8�I
���.K���	�ꞎ@..Zk�ւ�1�����Ԁ.�2��u,���F�$���������o�m�u�_�m.��c��M~�V�����$ݛR�nkԬD,u>��o��+�˓�\E&�L\���x�-�������޾q���=�Ԭ��J�1~
}f��/b��;�"*1���I��vŴ.c��z��
E�W`�u��@����r��c�X�����Hj<	�@cW�p��Hf��bv�N�B⢥��A0镖���B�3�܋�i�X�b(��C�a�#�%g���r��$|��m��(��_s�9i�L.`��N�awҥML������vNx����4�
���++�@Eq�yozQ�������"!+8:+_�,�����xӱF�n������d5�����t{)��"���F\2՛�D�zQ������bR��W����]�3-�޻�5��䟊V����3���������\O�=��~��
�!��17����{fjQ3z����$x4��:�l��ͼ�����-F.���E8)�Ծ��k��k�nl}���uυ���H�aL�+Ꮊe�e��7�a��C&�[�C��GT�q�����q��".;y�ћ��+��8j���]�D��:U[X�����=��&"�y��H׾S�6��� +�c�<���j����A҉���)��ei;��:����{<m�vK�Pf:?=��zNt�.SΤ��#��q1�����T��ѵӻk��<p����٨�8<��H OK:v��x���t���s��\Wu���I�-��l�]@�jȮ�Yߛk`�f�W	��W-���`��P+,�Ғ����H��z�)KD���p����b+-�|o,��������x������t2��_���0�d*��j���m�41a_�B��A�ꓒ��ۉ�ˀ�����=)����uUQC�T��w��˾.M��U�ӎv'�"��y��a�$�ko_(�:��v��R��F%ֻ��k��ׄ�������oȒ ��cٰ�bw@�;Ef�`k�'|L��vT�K4�n0��$I}�/AE��ΰ��mr�ӯ7�����w��Y1(m#�_e�d����5��d�2�R� ���b�-w6ķ�F��[�Β<��n��\+�D�EC#�u��DO���ʊϕTdN�%KF
9ш�������_R9x�S�g �a��a���6�D12����!��հ���Tr�@VϚ�����w�W�������"�w�+J�'�9y]����q����<�ːֳ�!��9;*�{�U;�� �F�o� 4B��%O�j�W��t���1ן�+���萸�+0P�=�1
����t�M��X5
xB��;�|ki����3����%A�-/��ql���H�����E�J���_87W��YI:0�n��ç�o��<�2��1��lrh7�T���w?����g,ɨ�|p�`��9!!����W����\���:K�&��'���ń}(�X�.���G�Z�\��G|��f@C#֠g�>��qZ���9m߰�/I�$��V��Ͽԉ��K�ma`a���F%F���y�u�6t����%�k�>	?҈pk�hZ��d��PE����)�s�RN{o��Y�T�aS/�ꖔy'�g����ۘ����D�c��R�!7�p��)��_U�y6�T%�7�
Jf�ROS�߯�# �0�E�E�RR�@w�j�&>�ԌP���,I������m��#��s���z�� ���Y�����)Jz|,��f���ͣ��y��)�\ ��HD�2�g�uV\���t�qN������L���2Y�O6�9qNC���3���.��o����_=�Ԗ�ʫ�q��E��hG��o�;�Y�$P#�g�O���#��ɠ{#���9KL������Y$W��ohP@E��I]t8�cn�9c�b�00ɢ���/N�������>5����yT�&�AbG�9�|K�g���{ԅiZ1uѴ1���s+�0����lR+��Xx�n��뼨u��KZ\L$L�k
{��M
��E�kOd��+-�i0�`�����7�eK�	)x�]0Ȅ
4GS�A��y��xrX�(�&��>��o���/�D37]��#���̯6�A�/�q��ڸ7�B>?��V@D;���a:S�� @ȇg��b	�C�2#�7�Xp�	����Ub4�N����Z�$uXQ���_��u/��Q�O�P~�됇�-99���-�����9���[~�$5�.���٩"��7P$�> �1���|�vr&�(v�,'ݒG/2�07#&���V(m=�B'X�oU0k1�`)p�]7��f҅9��63�wN.��Fʀ�$%�?�-p��d%~Q����:�^m����t�f�e������H��f��{����R�Ǥ��gz��j��qM�����
1V�A��H��k8�Ku��f�<�&� �����	|yw��&Ŷk��o�%-��[���t�O��b�TW��v�$ɪv���0NO�i�ڞ��/��p�?��/�mz�S����?��^�&�vII���%"��r�3�_����%�i��7�=o�d����~Yw��MK�H"3l���.m�v�ژDt�����m���a�\^f%�s�_�=Z6��`)��D���I�Y�*��.����r�")��	�j<t1�����{#�3��:\b,B�_V�1U�R���J�V�8�v%S^����T�Vω������#���J�n�M�����׸0,z��-��!��(����wߌҡ��f��"[��u*{l����E�E�2��E[,�pDv�bT�_<H!Ǡ�#O�-޿�!f��1c��|r�X�߰Wi%�,����1�^�*/nQz�vq,�67�L_�@��Zʟ��]{ؘ�|L��������g�j���&��g��{��<�3��G%�w�ƥ
Sjql�zf�t�*LəNY������ x�[{@��:p�pS�g�*�&Hҭ�{J�|�ػ��ȯ���T��lA	@��PN�U�[��Ԉ���4����G��f߭��S������E��:N�����h�+���3	�E���a���H�n�[�ע#N�Ӓ� ��s����3$P�0�Z Hޤ��I]}MN@��'5�H����M�C�,j,�(Uo\�{pͷ0���PK   R�?XeX�^Q3 P /   images/a8051118-2cec-4f18-9b89-ac75f15be4ed.pngܼuXT��6��PAP@�F� DJZr������AR�A�F�T:E���k�ffߋ��~������o��������<�{��׊2$D4D�Ⱦ�T��˓ti����h�-���sY�����q ����K-G���4WSo�q�z�j������	����inc�h��΄���4qC���A����ܒ֦��2L�puy*c��,�YZ4�������߱�${}I�߷��$�?K)+_2��,�LR�qtKxK��+k�C����Y���R�JtF��^
Bl*�β��{�+��>��N)5X�_��zT"��5B���x�2ˆ��E�	��Y}~�����;�/�=���ύ�l��/�Y�zJӰ��0�r�|-��x�$"�A���P�p|����Ƈ�.fY��xJd��q>�#�g���J�>�K�6$lGȗK��S0�'G�xT}�3a�7/teȸo����\�b [߳1$w�#08}'�;�"h�������
�ʴ^�����i���0��oaot��R	{3��Re�2(BqrIs����:I ��w���s/�7ѝ�P�gG���K�\�,#�m��O)�$R�WF����%eLv}�U��o��������M��������T/��RB��N�cG�ы/JV�P�þ$�̲N{{�N
�1��S������|����(/-�.%����WVJ�wdoU��<Ҿ(0;v�X�xK>B^�\���ƪ��\bPyiC����Ph�]h�����ЊM�?)����Q����1-~�%wUO�jE��r�7]��Y�)c�+����֠$�S%"���K?z���WhsH�Ȍ�9F0+j��Z$�,,,,[�@�;f��V̟^eފ~� \��](]���ߟ3d��s_/�.��eQ1^&�\VX��Y=�ⓘ;jg�"�ѥckWP\��#��d�}]N�]NZ���_����0����H[ZZ���K����MCMݰ�w�4�r�j�+sƦ�����?d�f���φ.�`�w$��kZ�.g1�	��x���k�0���&�dfa8<<'h����B�D �݆�$Nz�y�AXZZ:M�T�ʧ��:�=��8J�5�����������d� i��Ҥl̙e>1!!��FX[[;-?�}||�wz�?8ȯ�JA���U��,ܼ��Y�.:;�`��ߺ�% i;5ES߹��4�{߶3�PӾ��?9y��ںl���BOPJJ���ZҊ�5�W�<��f�9�����������6rss�MVL�m%�!Ō\�Q�����.q��\\���M���������ݩ��v@>��i�@�n6�fm���5EPk���{Z�q�e�H�;��C�Bm�0�헒�O����T�gw������z�A�&ah�`��Rf�H{�x���Gܻ���?��fF����㠠2U�^e�h�=��Bғ�HfG�����j8��˹mٗ�&~�ȹ��eo�=���0�5k�h�S1�f����G��?�)���j7x8�/���Y[�	2�tqToll�x	�΁��� �Y�:	əB�.���i���`�I�EE�F�d�3�B� ���tK4�f�R	�1+���2>� �� ���/i ߞ`xFjݗ��������_�眱A111����Ff�7�Pt�|bbw����;���;S�)�K
8���~�F�֕�*++=�APp$l���8���ɉ�������4���:�ќ�?���mt}���Y���[��/9d��ʕ+��J��7d3(������R�e����:��bP�u���^j��#��vr*����qv�	l�����X=W�poe��co�À�ޠ��bU3S�5�>�w�AWaX�S%���YF���3˪`+:�j@�C@���Ahۡ�7�F�b
�6HĨ�j�фuU���N��eȠ�N0ӠE55u����'��l�F��|��,�E��lio��?�l9���|�=o0�*�.�ٖ ����[M!���Ҝ����N�ڌz��ps��G���J����c�ӸP#������_$����F`�!\2�]�i��L�9u�'l�ޠ?���W@�0ñ%Ӣ�$N�$�%)�?j��ϯ��1(�r	�ɔ<E˽� �ˉXLf�W\̅;lCHK���)7S^�����s/z(c�l3�P]1A�]�mMMOt�Ѳ]P����r *��&_�0P=_�����j����HW9Ө8u����=��ɉ�@�<_�8�� ��թ[�Z�����*@c��C�vͣ����M�bZ�9J��l�1�L�fI?D)y����%UX�H �e����򆄄����N�lW�:�IHI��GA9���`����bq�~2&��E*  (a�D�辋BĨm�8�L�/�_����eZ��Z~��J͓�Wp4�@{���\�(`n�� �36=m6�B��5�0L��O�����.� �肪>�,���UOsD��� �Ν;cK�=���ݶf�L�X��Y�t~${J�$V89۲�_�d~�w}�M�9���>�S�_�N�4���U܉̎����_bѷZ�H�����پ�{������틫{Dݜ [�&Fm���x�5�Gm],�����7w�θ�!j&D-O�Z,�]�f{8C�k���J3�E���/���ӥ��,��luK�Hڋu�?�^���2�6Y��W��蚼m�31!И��]�C�bD��	q�%��dA��I�L�Rb=��k'�����5>{e��O���������:�~�#@��ѿӘk3ezz�':L�By�#��HW��z�΃�c}�A^?%�ۤ��t�Jr}*7�<
T�(7��e=�S�?tTU���9��${��0N��|��Ò�|���s��͉#$����Κc������M�p���S��*,��C�z��ߥ�/��j!��i����Ǔ�C^9�j�WX����E��;~x��}��ߣ�{��*E���Pu[϶��Y�Rת��)DS����J������ۥG���/u����6?�t�_:^M{{��p���Wå��M�*I5�O�P3̹Ub֗?���IO�{w}> �,(�N|��φ�h*+Z�&&0}=
��� {�������a�'�ʱ����Bs�_ 
�Ԉ�V>�Q�x��_'U�@@�
@
_���^%`�i8�W�x����ʇu�fp*J5�*��W�p%���N<5�BKG6�2f� P��8���n;�3b��_o��o��z��j?Y>��VK��߷ ��iJM�������Y��{g�S�;���kr��mfD�d�+��
f ��s���O\ �n�#�NX������eB�<	�ңH{�8�A��paX	hﻙ�����_��D��m��c3�B,��'� ]�۸DǍL��h��*�C�ff� ���\�Wv�D�AQߵk"�yǢ*�
�f�E���a�% ��V�`h����T1�x��H2G�*�X��p_��ʪ.�S}��s��	@�p�nU���B�jQ]��߭?H�?�6:S�hi�]�$�Ik�<�X�
y	���i9j)��C_7��J߱6Wͮ0�j� ���������`���l�R�:�x��I�`OZ��߽U#ܙǉ�է�S��U�5�E��eM�ƀ[��x��o�`��{�穅���CM�~�=�^�PU�p�6��OD���v��wb}�	C��n�&<NG���B�ߵ��R�s���N�Z�R9���1��WQ220�(������|̖t����|��K����>�c��{�F�A֛��͍�?�R��~9�-�JH`%#�0�) ��]�9Dp��u�^0��::_�Hf٨�yV
"������m[��&�(�S�5$U=�ބ�q�����&���.��̑�=4C�:����������U�-���şHHH�Jc�"p�n[AH���D�udG�v�����[�A	����ٰ<�~5�<�g��D��(L\��KIz���\�m�W���m��Z7<������m.%0\�&���f�m7bC��q�����	&qf>�4� �)���ܘ��`�l�r��4��?��'�g�VRb�:t|l�ԙ��6fNHn~��fz�dD����-����5�T#u�o*��&�0!��ɮҙ*���Pb&�F>|�$�L��R�a=�����g�&+�y�㋇�
�^FN^�Kf��m��G!OA�2x}�.��i w!��Q�Po�?꾘�QM=V�_���Ӯhld��FP��Ã1��C܂pt����΀3��f���'�A���x�����8q��F��u�__ z�_/�P��U�,K2E�F��Ñ<�-c�ޓw�g�T�%."0�Uk����	��&=�(���|���
0��5
r,� G@�`�����~��cM�F�iU��`V=s&q%��'0ſ�����[dl�r����I�7c�X�r��lQ�F`~q�H��vG��H!�4���v�p��v/Td%g�u�[�Fc�7��O���*�e>��N�JD���~\1����=@4oUM�����0���࿁@�YSS�k�C�OR�Xi���I��}�˨�<e�4��$۠��*Z�J��|Vu�0�ƪ�gKX��o�V-$��y<\H
	p)������/�\�~�;a�_���C�4K�����������w=��W r�tʆk��-�g�W�nn�M:tqدW��A8u�L����Խ[n" lV������imp/p�A�#'�1BŜ��"ėt���'Vh=�$����=�շ���6�G� �If��������B����@:�!2����f�eSAP&��o��<J����+�s1+�s�4��]��"W-PǶ�IQ�����j�)�a�| {N���sV��s�a4C$ڟ>�=^��h]R�2�`�1�q��l�*3e������>�����Nv��zPu�0&��R.�hӝ�d8��o�?;��b����qۏ���f�Fo�ܘ'k�FN>+���+�#�>�!6uE5	n�c����`Y7����P����q8�&q��&�ڀRa���q��%FH�궂S����$y�7-����r_���>۟����f��x��^��`����	+�Գ5S�X=�;�!+��<��\2ˋ�
Y�З^P�#;$��=��XBC�\]���mQ�TH/��:��{q���oܐ�YV�V ��YQt�";�E�
�3�H��O��2t%�2Қ
ʹG }�_�$v���[U�o�1�a���q{8S�YZ2�~�:�gY6fU���_�SmmmkJ%�y�	"�c_Pƛ$�:�����=��|0�oS�w��|�ag���uHI�2Q�zz
�����Y�_�,�l�6�Ku(��0��P�7��1:�JdlR��^�h�2\L����E�2@M���V��v��q˰��f�ɛ#H�7[�ŤM�j���Hdp(�� P�B|/�F�����G�U�q[a���P���/6��iC m	�� V}�#S��5�(����|��v��	K�oP���f9�`���,`�}�3���Ǉc�:��]O��Om2.���\(��mbuoU�\>r��E.����9H]�{��d���-��wl�w���|'��z0��,U�5%w./�' �y��ْ8JQ%�u�7F����x�Iv� ��2�{p�H�y�N1�Q���r���Hљ�MǕF�w��)V���@x����O���D��dV���eq� �P�FN(#�B�=��x���?��R�~�uɷ�<NS{��}��{S�5��h��;�.慉̲��mt�bᭂ�
�ҡj�#q�~�T��٩��>{�m(�s�g�%u�6���m«�ЏC (���h�{-�e�ݙ��m�^���:����?/U�x���L���^v�V�ԨWʧ-ʧ�R`�A��<�[��-�>hF���Μ���~>Z���j�V������&7PNKXl�C��¸���z��tm��2>B�J��H%��XyWn�H�>�%Pг'3x
"?�|b�\�K�t�666B���oՎ4ج�XVP��>R��Z�S�9A�� �_*�L��ܳSo�L(as�����zl[���xa�KA����xvws֭�B��h�74xw����~�/�w2B)]2��:��_r�>�L�Lh��Y\e)Ў������68���L �>P�<"""�YYYB�K阦��wg���ZF
qX\�iMQhJf���75o3�Xm�Ԧ����W�
�nm���i`�F9_
ؔͽ+k���~��n�%%x|@�mi��h�������5_��ĹS��F�d9���?�v!q��1˖�t�G0!���k�2�o�C\Sy�ُ�\L;�Gf�?��\p}�Ԛ�ڊ�z�߸���m 4|}�-���
�=���<
u��:u��#q��qr��g̪?��>�Yh+Uk�=䬙���;��!$��*󖷷7�V�IlW���S�&�?����9��P���>����F��@ߖ/m��sR)����,6�����z��<��/�r�Y(u�_e�\�B���6]���L%1�u�:=̲���A���Wv��
l��W+���"��{�ng�H��8��~�r���{��f�Л��d��jnmRn��qv�k+S����3S�b�pϢp#�@�6�4H^qgb�vr��@ir��< l}vK����_��������H�G�]�4l8�/ě�z�ZTд�q��p�	�P��Ձ���6��K_���aTú�hλ�þ;6��{n亲Ce*Y�"o��"�|�B�?�����|�2���?$8X��9� :�4L�[uE�7�{:O�z�� ��\ڰR{�V� >�J���4�[���J;a�l.��O���������"`W��b�)ٳ@f��+�9�\��n��Y>h���F�}��~V��dV��� m?E��Ρ���^�A�Q��уuacY[�ŁG�ɴ0�5����xS/�=s2���/�tz��W�c>m}�g�j7�(
WU (1,bF�+ ���$@߄ۍy�c���e�ض�u�\�R+<{��8�� ��$.3��)ꯞ�Qn�7�<&Tٸ-�`�<҉�������R@�MM��Nt�豢���Z_��	��8��t�ڄʄ0��7pѻυ�INLW_o��m^L"\�V/�:i�-Ӷ_�>BCq�{Ѿps���d�[O�Y�=x�V&�S�I��Qӻt�0q�iS9`��U.'���d���*�л
��\%�G����٨f:V:J�)}�ti� r=�j��Pc�îN�Z����?(	�9z?3XG�{�c`����GԴݸ'�Q�,�p �o���@ wȢd�
����wj6��<��]�:XP���(�n{d��l_{WMNF6���Ը9��
Z��j����!�>�[QU��[��}7�ϩ��BI��9�-����������@�������KJ�����e�x<����DkC:��?�V������ ���3��ס����e|�\�4�3EӅ�5�MO�FPA��|Xұ*�O��\ǩ'Ƅ9�R<Vr���Ubu.>M����V=����)1�h_ܡ����5��s#ӏc����j8c��U(����+�R��p��S���E���I��9sn5�Lg⥣�)gu��=�ӿ����8f��x#RI�ķG������%�	$�n��2������B��;��޹JФ���v:��� #��ӳd� �vHQ�ޞ�T��o�t�F"Ľzur��7R1`�ÍW����b7�g�t�=�Z����=����VT�BU�ש{7s��|(9�db�US��2p� ��mܞoG.��
rsߜ9l��D�^��)D>��� ,-��)��-k��n�ii�)~�{�G��	 �q����J$��ݟ#37[؋�W��T'���q���l�Ƿ����'Pa�r�	�	�����`wEm��O`���(v�V6�B
��ON��]-?�m	��Iݶv҃�1R��Pۀ�:!T���;�}$#R6t��0�
FYhqUU�����d	���Q�6�y%]����)·��ч�7č����V/$X��A?�XD��|S�N�?�* �z�%�&��k9�n���3<\��mA	x^8��^DPq�؜&fo��ӝ�
?x�:�\3P:����nn���?4߅�?���͍zn
��TZ�;yu����9�͎)(�D����H�V�v�.�s��W�5ώ� b��6neQ����? F��嘇`Ӯ% fc����ۿ^lu㰩����@��} ]!WR�(����$6�eSw���_�P�Lp�0L������@bHJJJ�cܺ�X5s� x�>6갍!E�c��K5��f�>u�ڗ}{4:bц��/�I0��N5/�Yv���.�R��g"�^k��9W,����1˙��
kk��Y���Q"�F���kڃ�E8H�������p���W@��&��I%�.� j��;~��Mݮ��٫,��ۣ����!af��X�>�X%��9��p<�80YA��JЃg3W�'��M��b�?3��wV"�GK���˿3퇵L[����8� ���)�<��,Z&[f��n}̟���/N��	u߂�'������63~�hKHG�2���S/Y`b�உ�/$��`Ad���G���_��d�Dk[�#��wu���/��8-?�r��n�ќ�q�Tl��U �b4@�:�������K��������&�^|�����@�ok�0#�����јu�i�6(�Q�;�'��Cx[��V� �������,�����0| �V�04zw~����&T%��tˮy�I��0{1���WF�+�%���m&��s�W]��b�7_v���a�Me8�^��*VYc����x�r����4��C�)y�+i�Z�]?��6z��u��xn��M���r�d�R#�FN��/���������-5���4�WA|	w6���,����5�W��כ�����������]
��	�W�,N�lC�Q��y8����?���W��/��|@��B�_�~]Z]�����$9�~Ҭ�����Y�4��B~2�[~�i��ځ0c�|�5�u2�,R"��~ �ב�q�����.)LQ]���&�������Ęo��m5�)�r1��*/6=�i ����{a��כ�;=��3c�)nx�0W��?2�g�,��%��g�w⟷t�5_�^�[M����+�\��c jD��P�k�<5`�&q�*d�е��?1!ZD��{�^�m�������K��L�O �[C�}}{���y`
�c�8>�|��ў�\	�[jg�"uF��+	�qN��m.����ړ�:̿��]�J�����we�SSt����aͲ?퉅��O������`�y�����n̈��T<����cȧZ����kJ[9�ɸv�{�	z���q,3\��¶���~)��xӔ;/^�P�&���A�ҳ�YJ1n����4޽��)1��u�:5��0��fC�Q-�_�^�
��ik�/J�ݩ�mm������4�M����ύ����}����jg�fm��N�A��e�߀���<	�,��U$W��+q�v�إ�%����|(G����Ϩ19�ӵ�T�>��x�t���b���>�i�H%�Kj�T1���mWL�n���V��-�DpO���&��J0�m��X���]�f2��U\`r��vW�[��+JhE��!��a�-��J%���Q]@I-�����4���]\�.��Q��g�#�PLBB�HW������>g��wB#����]��N�l��I����vi���O���T��M!/Qa�Чò��I�"��|{��� o�T[�jQ_���z� NW]���b�=i3����O�++��{�i{3ƀ�<����:޳��[tln�]�|'�/���Y㦂�?��H��a�,˛	��ZS#���ɔ�VS���ޡG�G�YCz��yE����!n�S��.cx7��ǋ7]k�-W�gg���?���I�=�	���F���f�6�+���M�y8�d����0x;
8`5&�w)v��6���AF����c�zW�;|��NɧZ�43��.����htJEMG���aQ,)n����� ���ݕ�<9���r�??lkjj�2�E�;v<t���|�:M�]a�}��k�dejj<�j�����星�d��3�QFb��HJJ��EK�U�_G��S�u�j�>#�Z���]��?lC�s�s�E�kބ��Ol��������)zS��kj�RZ�a�z���ԁ+�P��#��N�O�K�� Ԉ���=��y��n���RR�9��8nKU	F�������ό�a�������"�gn�t.KQ1��E�+y�+y��wP^Q!Z�@��#�Ȉ���/�I���2�}����ws�
%x�88���oS��2����@b�	G|��#�#������C��u%q���q�� ���/?��}#�K��W�I�`�j5�k�M��,|�p��:�!33HKK���j]5u��KB/OS� ��?z�#<X#�v�����[�\�wһb2�5�
1��/�6:�Z�7�ٲ�n�t0��x�X��{��4���D�%��H�:��0qa���7û2G٠�?�p���A78\ [B�ҵ����-��l��m�{�T|�W�0�=�~p+=3�Dwնao>��O�������qBLzUؙjt `@4���&1�$�����Ӓ��e:�{m~�b0�XR�~�@P_v]����h[��X[�h���x�"��E��������r�K��W'���[��+�w��˿7PI���U�<>��'���zJ����|z���ǝ��$E�R�qK<V�VG��|)�_S�V��Yd��7�>q6��ޒ�Z1LQ�Q�HeHG0�ok
6n�P��%��Uc��L|�q <����O�av
��蟄�t.XoA���'.�ʒU�Y�}{�߸_A�#����d��v���<r;�����R�(��p3�F��_������D/+�8��e -�i�����09�#sp�r��X�4�{�2ix:���1
{�Μ�HG ���G�M��p2���0�iYՌ�I��{I0�/��|���/E��,�U��~���v�������n"ѵ��q#O�	"��N���/ �|@��h}}���h�L~��|4�s���ac;ZLe@�X	V?�}K����)��|�������8>�FP);�P�1��z�9y{˂2�*hJtv �$��녪�E�B�.���on*`N闏W����$<>0����[U��� �<j|�U�S�͓  @�3x�#ߞ�)��g��/�K���쪇-���?��4"&O (��朙����cύ��k�r4����"?�bBC�0NlW��Xߋ&V�;::�lgtX��KmEt�6�j �q�A��cb�M,�!E��%ymw�X��@�� ��Tu&��g�������~\)�w2���Q=����`��A�,��SO��c9�r�|��X	lT�����z�?��M%����� �:9;K�ȴU� �w��xS��,��ɑX����زpz�*i\'8����f��^���@=§&��>�i�2޿A4,���@׀Պ��,4Ϣ�c���&P�)���_1��gZ�W9�z4��&%��]�2��/���l����]���~*������5�����.���1}'{+���E5�։7�Opz\�aɛ^	Bj2���Sa��"���B���3^������_�R�\���E�'J��D���j�-�p��b�^Wy����>ʊ]�'X4RS�=S%W�ܲ/���/�_2�W�nU�#��AxC�Mx~q�!LD�JA_�������FrB��l�a�"�9����<�|���� ���P�ܚ#�KC_��pA��A�V�{+C���u��W\�����N�p`��C\�Q��!�xN9wڵ߃b����Do,t�í"����z�>Xm;���I^nn������p������E���,Zcw!v���o�?�D�%�Qg�L�,5�B�l4��IB�.���.���Ne��7=�As��9��"cZ�I�/��@�����)���Щa��hO�I�d��dy�������j�Nciz�������fS�:���<*��(�rn����{n�Ƽ����2a���_,�N���:�eX���t;�gWAl~Ğ6G?�?(�֮�S�^�m��=r��Iti��;F�1 B��gD$u�f��'�Bb�꧰.��L�=�_�i��AO+Y'�N	9����g��(\ٕ��
�\(��O6"�=3�%���~�1o�F���`���9��D��R��@e��-� ~�-�D3S�w4TX��:|b�O١m���@���+JfN�.��3�&��|�)�C��������yc<Xj~q�v�'�U�Қ��UV��N���"�2J�{Q?�~[�/[=�˧ڽ���-��Bq2^�^]׬f�=:���Ǽ��=�w\��ݭ>�WOj��e��|Q��l�@�l ��\���<Z�9*m�-ٱd�8��X~6�Ƣ�ѳ��0=u4� ���ݎ�ŉ���5lo���t�z�h��W�4R�F,$�)���y���ٰ�"~�; <� A_޸5L�֊���U?G���`��1��T�]|�y�?���=�C��S8����}�ɕ�K�|��)?�b��{�rb�{G�yH���C)����y���a�4f�$#�S��KC���p�^D�mS����e//s�:�ܩ��5�:ݦ*��t,��t��k̟��p~��Z-��h�x
�����)�f��X������d7���k�ع�tF���;�^���`h�9s��\(f)����;Q V�$N�%�4��_�E[�q_W��]L��/���L\p{�5n/�^ �����;�7��Eڛ �̎��=�NQw�}׻2��n���ӭ�5Rz��v-�k���/���n�t�)!���k�E�`=�K�t�2�՝�d<���Yt�pW�]��^ER^�;n��K�S:�ήY4��T<꼟^��a�����i�1Buz�B�)^۲@Ț����M�Z}8�Yx��ɤ"���26Snp�U���Ψ�w1w9�t5q偂t���ܿ���c�ާ��J�z��n�s8Qi_u�S���P_��q
��^��Y���A�a�
f�|��-}s;H�g���:��R]Ԓ��~�����V�+6\{�\2����"�"�u�ٺ��9�_Q71�������;Jl��w})���Y6B�re��(NR3�u�AL�D�����V,�56�t'�-�k{��1�@�,�Q>j���ӣ"+�6:ץƓG.p���6L����	��/Sa���p�N
�����T�LP�k��-����	��Q RG��[����<���í]>��7��$O&���&z�.����h�>�Ҋވ����!<wshxx�ݰ�]��Œ���z���VQǏ6G~��YՕ�ke���O�&�5���=�0{��(v��C�ް�������-<[=u��@��S��M���+��4j���,֞wQ��������o��:j��o��h���v�?R�md���ԝ�Ezg���3�;`��x9����2p��ꢼ�_�M"��VNC�������db�r��C�:�{������g|�CѺ�ݢ�J�YMT�9d̴?�<*,���3��Ek��?�e��ssr^�Ѩa����4iߖ[\l����HE���;vz�K��j&W1z��?3p��[�6ޕi���L��̶"4��=�����trZs�ӱP��FR�Uا�TW�,���Z�ƄN���G/����1�k���|��Q���¦Qv��3��ț[D�X�CN-��@ܺO,q\,������ɂ �F�|�� 	�t����ٻ,��B�l0�R7�UJ�x��8lfѕ�
�:Ql�%�FZ��O	;Y+�Ш��v�8��X]������gĔs��}� I�t~ecC 
Nt��VL^~>e���2�����"曗���x02�nB��X'�>��{.�m+�ώ���8'���*��'���[&�(JH}�Տ(7ZX���ω������{�InV����W���������ԼH�哖4$��;I3�.5�7Yo��`�׳ 2�+]\����)�$� �
u�{
��k�}���QG���q0� s��͛���R�Ò�2�^����*�pC�l�$:��mӰ��GR��E���][�Ṿ^!=�ᾆ�� �Փ���������D�����N���J�#FqM^�2'�K?R�U&� �������ͥ�3���U��%�z���YIg����z��I� D|��9�!�79�h�����V�!|��k`z�0�-}|\[+��p�������6�I�5�{�Зϯ��FŌZs����қr��[7�7��䢖��<���{5n߷�'g�!�#�/S�~yb9|���7����7�ḯ��� �Tἆ���'�h�?���Ү����J�IP��8D6�������_� D�&�/�7&ne��"^Q�zw�A�����å���n22\[�=0Sܛ��z<1S�vn|�������{3~�﫫�W�<eI���
��S�_a{��	U�@D��D?f����.�����ܟ�,�G	?�R�ם ��g�iiV�g5����n��kh�������Ό���F~g
=o{���|C����c����x�3�
|���gˆ��ն�~��4b���sŅ�O5,G���e}���+7 bl��b@�t
�ݥj���y�U�W�1r%2�m�٬���u�,!�ت9�ea��7�i	�
�I�����X������s��>onf���S�6:���;O�;<�7U�׬�]�ߙo6<���71>Z��>�������ί��p��J�r��]L�2Sܨ�Z=_M=��f��X��w6S�w�D�zΫ�<�L7B�D���i�/泌�E
�}0[:;g����wwR�\���0�~�ȫCI���.�u��Wf�ǅ#��^*�^�~=�q��dR�0}.�/.�����_6��|�~�-�0�Щ���� ��X5�p8���D��L�,�1*������^;�-��������Y��+���k�}͚q�����p�_���uRhac�_#Nu�����.F/UT�괳�#��X�/��!8�`�Qs���X�h��|�~���?�4,utt���j�J՜���{RUD�� 8��e�=����պk4=,�mn�xn�~b���h�+I�c���*S�H��8�e���_�.�#���B��	�vr�����c�D����'��.�;wמyJ_3����
n�0��H���tA�?f�a32�w<ni[GI}&d��/��mD)r��*�xwO�=ڃ�H��1rHz`�6 �m"����06��e�l71?�D��x���I���M::" ��8S�=�;2j9�QΉ�'�׸bc�߿u����ק����坧8�yX��֖���*{�l������ݴ��!"�nۢ�<$�r�&�l�{8�E�E���q߱���0|�����R��R��x�j.�9m˂`���p=͎뭋PP���u����ml�l��w@M�a2����I:��o����������6�$O���}!f���Q���f�ZV����i���^;�����3�������ć��`�W*!���%���$ϡ�:��V��;Y�� ��:6'�A6�7�������<�� �E=rDmU�j���������1�C?�b}��Z)� ��&����\�9����6@��h�9҇~u͛x<N���	��?���!�G�e�"r���@fp��=�MYt��5ݎ�'f�ƭ��p�9!�H��_T䆸��F�C#<t�������*�;i���E<�s�{��c���Lf#y
�KR�?6�VL���(���GLb�3B�,�Z�R/���<�������i�U�s���� Ex�jvu��[ی�U���c?E1��I�IȱmM��$d0��\1>w�x>�7^�qtuZ�2�-C�n�y��EYs�H��~�H����Z�v���>�õ���,W�Ԕ���X2�-�q¤V�Q����X��,��+3���~\��������>�����iRL�`
���c�we���K;�S�9_�F��槥1�W|�|.�X�Q4���f{_��!.�v��ɣ$r�5+�i�ٱ���|�-��ȉ��!��?�a�	��WV
<���`�K���&�{�1�����/�Z����t����V�w��G�U�8�S�\�ޟ�b��B��9�yp�r�D����:�]Y��'���	d~+��9�L:Q '(j�D
O3�/F�}�|<>��Q�\X���)Y=f��ҿ�*W���"���ى��܆��EX�>���3�������5��->���iJ�7U%��u^��ع���υ����;2Q���_�oω��睝�D~�ډ��[�{K��NnmTĮ���ky��_��N�.U�����J����2p}�(PF�S��u��wY.|&�������Bt������ڞ�C�25�J�1�k洔R�L/��z�=1�Ʋ�l�Qi�c�ޥ���m(�LXs�ٿ|Vy��c9 ~-��;VL��|���{�
�(�$4p	���؛rZfe�WN*��mp�91�
N���1���Hvv���Q�Ī"���uuC���蹡�B�X�5QsG@�MMM��45���щV[�� Ԫ���z�>��,���=�{#??�2̒��{�V�Cێ�t��"Y'y�)6���f1A�%�H�lšV��!=��`�� ��
W��]]]�3k�'@�j�Hy�$k��%$&VXOT��++����$���X��KE�G�F"}P-@f���`�S��ߩ����v����"D��y�����%�O�z��-����oQ=>�3����p^ը��
;�t��v���R32J�ݪ��BB+�z;h}����}�����v���*�ja�3�Xq=x�>-"��ǔS��d���F�pbdE.		��8*e��uͫ =�E������R��������[��?岖#ES�[�Ï�Ó���/�r=yg��A��/n�~FH�1�\��J:�.Q�$:`�Oq�IeeVJ����֮J�1����[1u�)б�ΐ����R�N��v��BW�D�f�j?�u��D��Qkp���,������\�zk���	O[\�{���3��YB�//��ūf���U�tE0K�+"��ttt��b�=Iª


�S�O���_i��)dS�3ɱJY��$琕��8F*�:8Vv���	���-�ؒy̌��~����_��?r��������~��*)������_�B��O���<�i�)E����`��3CL������,��o4�i������?v5NN��L�م}�8�h�ř�]���
�Jcӗ�w���T���+�����h~b���)0��a�g�L�&as5�1�Ǐ�x�Jlqsnj��DEs
#�j���.+M@ �G3���������[?BJ0��]ؑ���+#��*	��o�q2� �%���,����h�z�G�ut��oJ�![�G+��u	����������cK|�BN�A��HX�m'��&HɈ�)�h+p%��a�ӥ3����Hu�V��Dǚ�K� 5���6?�~I=�)7%�^)z��� 7Eq�}��t�vss�v���g�\� q&�ۀH��Ҍ����7S2ҽ6u���d��lB�m-b���>�������7��'=rڏz��x��M����y�G��iȀ�z�3��!�=��m��+���t�o��?{�_��J��jj��8�������cg?7Jb���=1H�P�p�s��3R�M�']+�� (wEb�p��G��Zߝ���l���^��� (t�6�prP��ѸW������}�p�(4�O�|��"m|b����ܲ2���r˞,�.��FF��x��ZR˽��59	il\1������{��q<��hm�y�~�U~�����+��o�+�;%��i �PU�hT���Ff�p���:4�6R�m�&1���=��b��J�v��ž�hYY�D�I	��q�R^�خ��_��S��&����w�>&&u&�Ng{�S9ޕuΛ�+�%��$�ŒN������K�}�U�2�}�iW�����Fw=@�����ϕ��9Ǵs��7����O�RZͯq�*��D)��`�44O�&בxdj������w�^A�|�xA��1z��u��g��0Ѝj�[Ю��6��~�3;z2��$�!��������K7�g��"++�����H�r�s�;0X����6a�{��F�C��49,�_yͫ�h�(�r]'�������_R��������T��*�����]���ž���*���3���S��0]����"^q�)�y���IA�I����W�LV'���-*q��&4�.� ���8r�W����^0
��'_/\��x�<����ǅ��س)
}���ZSY�يk��y��Kv�\� n�Ȯ4a���f*�=�}-r�s�I�$'/��Hٴ����1B�ܬq���(Sm41w@:�h���9 J{^@�[b�CCh�t����g'����.��&1K����?1���&�;g���ҍ�^���諫��1��x�F�4,�N$�>�f4�5R`��䇵�}�Z-E`�婎-�V[�7�َ6��'|t��sm΂xVWU�}������mU/���}�v�zAF{�,W-4&L���,3ROTL�eM?���5)��lݟx��N�6���ғR��B[{��m�EP�D$6_E>r���6�N{U�3ZR�� �Z�ՁgN$��u�-��g\�y�c�{u
b�lt���Z�T�\�$��Wu���C�K�� 3����I��a�섕y��QP�����4�y!���'#��L�W�j��s#�s"j�0���͕����ꑂ��Nj�qc*L�#�r*
\��.���	_N�A�F�+~3y6ĩ�9�Yڧ
��祥=����O(�䰯��!Y��rU���N<�["2g��|�>����֝ �ݧ�\�wg}��S@�Hn�P��7�D��=��Y�/���|\>L�gk�Kn�lJ���o��ҟR��-2��V\RRbck+�D���,2�-��L�k3��xKSu��r��.�t�BR�r^�O�1F��@���Q��c��[Hs@s�D�H�<���\��5͔���z̰���f�[�����C]�H�>|H�v�o$9ǔߛ�z��x&��ȨmRk�b�,�ݤ�3/��W�>	�R �u;�>�F��V�w"h�BH���.���Z���}�`��kc������AQ���4���>��R�vI�}�����E�J[����ą��>����r�n`�����J5�t�:����H�� �('c2��b��DԽ�p�����EB�>Q[�'��w<�I��w>����)wA����P �\���#��ge���$��Y)B����5@jd��Ƴ�D� P\.��'�s'x��Y�6�)m5��bL�F�=?\����o{�����'D �kIOI�� F�Ywҿ���:����W��W� �<��2��-�;
��Z*��nw~�ސ��wn\
�����=�K�>Є`Zo =�ҝ�j��%��x)���w�k�9�O*����@�c�)*�r�����H�����䗖/:E��P�V��?��k6qsy�imnT�o��j)�f�7(��f���[��o �#� ?�|��k�u����F7��{��S���L����z�Eϰ�.laa1����#u�T��!s����l��O3��]0/]\V��#�t������n��o��H64.X�B�*�B���$��U^����O�)	xNZv���c`��f���s�A�k��&l�%J����������;]�C �?(nw�c~.W�%�\ް�t�iqG�*�fl�]��}��s�{w��dd�j8T�±f��"��pw���w3����l�֚5�	�����ø�9<���e3�����X�=>�y�ʤ����UxBބMsK4[J(S������ͩW:P�e��F(���:��u�h����;>�X6&��3��4�C��F�%j��<i�Eŏhu��_��o,���Շ����JQtj$mD� ��[b�T|5��N7�!3�O<�����x{�Rv���(h��V�S?�-���1M{��	s <�RY�۵� �wL���u���d{��y��^��I��󅀷��ɋ�+��	w�T���<=�ő���(sak��C>;ukN	c�[T�\/G���`����4�}�S����4R�7��$��w�R72��1N��=:ʷ��:���W^{n�YTC���^�ύ����(���u�Zu��~����rj�R����U��-�o7X���U`��ҟtj/�`���+��{���3_$[\[Ӈ����Hx�K�_ӹX�W�9y��w0�e����x�!���Ա�9�6�5F(?J�_]�T�e#̨���?�(�~�JI)��N30���@���js�F�l��i�,�6��<!�r�ÈJ:u��ת�������^�H@D��D��)�����,(J�����X�gгrm����VE }�q;yp]i�{8+���ϾG��,nTY�n��ƃ��=�w����Rf�]<���¤2u�m�^��`\�2����+W2E�%�Y�QD�ST�;�*��V��O	���U�p��Iy�^��6�Y�Pj�l�W���!���Bf-��ʱ��G�4I��?��ܪdV�=^RSz^�]Q&�[Yko� ��D�sǋ�X��n�����;ݨ��}�D�Dy���?��T=��w�O�5�Z�Δ`��J�R��HF-��{�nDg�O�ц{����G$p�2,�!��f@�58 ���ۊXrN�s҇�V�@Hz�����e[>�e6�Ċa�me��G��T-�����6�X_Y�9^C��ܑ�i�.����1��G�Jk��ʷ��H�.+iƅ��˼�"�ҫb[��Íb��W����E<�|U��J�ޝEk��T����./?uw�x��� d?C܃'����t%߿�gg8�^�Z� ��.�8�� ��"~�=��BBT�}����|���
��Tⶔ��<�v$��4�;A�;F�Eؔ


��ZH\M���u;v6{�&7�3W��#�O40��o+RsX�j�z�h�E���h�*йsp��mpW_�f9���B�.%�Ig��
�	g����F<�
���}�q{zn�����Ts�,3S@�m�[�"��2���_���B���δ6�|��=�D���3I��`�e��6Ov�aO�9q���� gu���6�,����cb���p:����+>'{ɞ��bL7Xd���@����i#n���%z׳��������ӱ��qVj���RW��7��҉�V���|Ǧ�ig+�^$qA�����,G7���*�Mt�yG�2_�J�9K�(]�Ý�ҡ�>�Ƃ=n�q�)������zc eT�� ��^��W��[J��Ð�+�~�Y��J��;�~=8�w�М�1���;���~�>��S7D���v�g'���h��{a��������a��_6I��u&G=jRD1�����x1G�ɡ�7E���s�"Ld��[�Ȍ�m��>�S��TM	����=\*�8���S��sI7��YQ�J����
�`S��iE��p�¸F�����j�$��="#,�8�^L��	XG����}#��������@�Z���9T"`�:\�?�|�ɉ��x�����>!ynS��B���G.�.�z���%%�>��Hŋ�#����-�yV]�\��yUU����M/�q���6�����>��Sh�0���|/\b�`�'��
�{�"�wO�;�OCr��I�/˧��+������)�X[GNS5�\��5�q}x+
Ͳ�ivC*��j�X���NF�G�?�B#-y��ؕ��:�o�f:���|L��axކ�nVi�G`�"��	_���Qb����<9:$��l^��4�C�p�����`�}BxXŏ]�z��L@�5��x�f#�.xV�5\�ah�L1�̘��\�v�V�t�3~C�@py>��y��4}w��V�?SV�� ��s��@��U�p�&�jE��k-��o��]�[?n ���3�U��RY�ۧcm.�M�6ֹBLf��eI��{<��-��xC��AT�w<��١��e�CN�<+�8V��V�S��Nr����b������E ��e��qս�b�gN|���~�����f~�!���Ꙑ��}ѭ��{��G��r���� }�;ו��R؄�����ɭ�Ï����	Z�j�^��O��?��EtӾQ�`S[�PD����|t�o_��(�Q�~�`5�G��4 b���(�#�Krz,oR$9��Al�����%�]�Ql��{�Yݷ�l�(�L-.www�SeX7L����,Z\4}'�u=IP�z��QΌ�e���U*�:VI��!���mlM'���5b �*�J =��~��>4~#[MeD�pK/�w�: NQ��[ޠU%O�:����U��y���<mp���-�OȤ�H;��~m����Q���Y��������Y>�8b�����P��s>K��Jb�.�k��Ϲs&�v����_�;o����Zců�:Di��[���.�bٻ��1Y����?�N�ݛ�yj����y�9�bVcSV�����-[���B(�����E	�{�!tI��}��˶h�O��(yk������zn>q^�"����?7�n�Hm��E0ZL�eփ\��6C�U?�6��Ye|(�y���O���$HKNNd�f0�؟T3�:\����|��a�E��9dNZ>�v-�(,��V�{/�2,��Sγ��i��ï�T�+��K]ҒF{��м�u�>�8�Re������I!�2�\A�ǋ�$ �v��f��ȶ�����g��q��\y��a _�w	Q��[=��U-�WJ)����Q���GN�ݘ�h�j:�H�FeX�q�1|����C�o񟆏33�yb�)Û�k��q5�ZO:��NL����� �th�� 7ǿog�90���h��f�r��|�'��DD����=�����e5��=,*�-�~�� m���^Hl~�	�1����Ev�$��#��kk^ù~�5��ت$�S)dRB�㑾>s�b	]���dTZ��	:�N6\��ڢ��I�G���AM��]Wm�<�K�s ��2 r<� �c���n�7?ʼT��c�M�ӿ��[:�q�7���L�٘�8��g�K���J�����
�X۸�S{ԏ[H����PYA(�=d��ؗ0�e7�(E�������v4�VZ�O�u)[/<*��|g�5���V�^1�q���g�� `�sAѰ�כ�kR��d���1=}H>oK�P�ۛ��ss�U9���_�KG�'v]��ܕ�QRW,�����DP �~i��]+�X�Li��`c����/涩(<��͌�"����ޥ� ����>*�؃($��?��E��H�6�*J�m��i�W�}.�+��K��Xq�*�Ap�x�,�e��th���&�Z�6�꯽�n ��Z*m�Vs��qsТ�3&|���d�'�@�����W��]]���םdƟ���;�����Ԅws�~��W�<��XF/=9g�ԖQT��ϫ$8�I�4�����7��<��ʭ�p���B�]�N�ə���0&#11��svJ׫�bf��vV�1�~t��%�G��9�{g}C��S�vVKQ���H"�{Z�=�`�.������#^)G�,�(5f��M�� �M����C�ҧфӻUlR+��5���=[�c��-%$2��s�>,�s[�� ��Ɨ.��������^��&��]ثA�^���ԩ��ݥ��m�,P����W����7 �5?Zz���ֺ�y+-��P͝||����Z��U�fΣ�G�55�M�I���c�M�$���x�w�R&�FY˵�%�n [$���"c�����1T��9XF��x�;r��-�����ک` ��q���?~i��.����6K$:��S�����ƞ��g?�@�\L͛I�ŷ���mk�X�k�~������H�V�_(:lXN�ם�&���U-��%RJ@ KZ2;����H�7��n�t�O�6+�X{����0��p#x��㲫>kmӶ'����̪��ri(������y���/��*'��_��Ns���u#_d�	�&��!��h�&j�[���2��X������.��jj@�&i�J�o�4���⦃�9���ҙ�dY�<���}�������u�x�M#N���h��Ĥ�il��U���v��l���4S�ˡ���8SP]�9�tS�����T�)�l���)��,�WĲw*�-g\̆\Y��v�	�S�|�걒�apB��"#6�0���`!ya���&��^9�o9w��:�3��o[�)��VPvjl�
�m�;e�]~t��~�
�I�&٦4�).��Δ�����8ǘ�0�s� 5E{*ɼK÷�k�qG�+'�j�Y:X���ouɴ!(�~Fj�>񾷠ڇ���y[��g������~wδ�u�HXѪ���;:܎16�h7�� g��x.��K.�Aұ&g�R���1
�2YH�
W06[��t�����yLIG��\5Β�����}E����􌥌�ؗc�HbJc�p[��!;��8���);9���3��6F���&	O0M.�ćVVU��$z���s��8��᰻��\�r�@^�s���gZ\PU�tGP	&�������� �7CY�h?�Y�q�0�$|��.�3��2�|#,
��;���#+<�	W)�[Be.3%C��%�;('��=H6��|�S׷�z�gjbCB�ӞL���Ís~E���`i����>r�����#V�K�{�\�<�p�v]�0�\B��~�rIٝ�ķ�F�-�o����у��¥��q+ޡdڧ:��	����#�U����1�k3�+����o^�yƍ�����u#�O2Ϟ�%.]��lr^�8y2%s'7��i���l-.�s��>a�9{o���$$|D9�e�آ��Ҍ� ��
Rqƨ�%��!�?:ZHݭ��!�;��1D��aIפ�,�!ޠ�g�]�N=e g\��Tr7���3�W�����W���n�+�����sO¦��R|���Oa����;�Q}=� �}����] ����z��!ʿ(WFR��,�9��ׇDOԌ��)I�'���\�_�+S����Z8��4���ʡ��	�z���v�_��Uh	���!�Pf��	-F�Y��n"���XV�M������PK�`�=��I��&�� �����7���ȁ�n�$b""�zל����Ӝ�72湫Xφ�?��b���;���
B{�dh�7��)����w�����%#��E5���w��<�#����Ӽ�oj�g���n�?P���Y9�dǼ�6,�Y��`Y��#�f��I.B+�/���l��ws��5�= ��}��$K�<=_�pl��!B�U���*���rs=��O�ꛞ'S�EE���CEQ�@�q��������I��Ȕn�3�|�_�˱~'\����Dgh��V�y�x"�#�П`kJC���E�����v�vT���/}��D�J����K%9̙*y`ض�z�RF||U��V�'���b�"o�`�}��L�V,l�n�}k�{�9q�Q�rެ��tp)`�e4*��?1�S&@�hژm���X�rK\TQ�;�a�86�Cn;�����i�8ǌ��٩?r�`[�L����2X�ZW�3��A����(e�Zu��g����2���\T  ����o��5�߫S�  ���_&Ѳ�?�Z^��9n1���A�����5@L��_p��nD\�q =+��)��͹��qy;ή���a�,Iy����1n���j����}(�Ӯ��2�Fe���n�ݼ���>�"ͪ0������s���Y�f��O��)�0�Ǫ�e3��"K�!���Ty��qp>�v�I�un3���_��q���͑��"���iP�{ǌK׍�������t{�r�`ܫ:C	�j!�>[;��_�����7{����Ja����wnζ����ݹ>��|��J9��S�0Q��)�Љ��x�vv.����W�H�`qd���Cu5�V�.����d��M�2}6��	�& "E�S����^ohu��%��X�J����d�6�K�h�[i<&��|\�4u�!Lbe�URWD'.sE���=O}S�W�#��'�{���r��x��G��B�����oｽs�n���a��DV��A�[O�������qq/\-W7Ma�T��&���r����_Q�	�hs��������j\�}��ɱCm� Y��J��.ehu�p)��ы� -�������N�ȑf�a�y�?�ܱ�Ξ{б��!��r�ڮ������/]�cu�1��)W����$҇nT����4գE��]�~�O d��}�g��{Q�^~��K���@���"i	�@zf��\�������b~�Z-~d�o�r��?,B���Z@ aϺf�P����n�	��o��<ݼJ0PW�!}d�M=�')�4X�r����6ozj��3���Jk��>��r�̓{�j2���ʍ�O�^�������.�7�Ԛ:rT��_��kG�<����؆��!XN
��s�7DK��z���:?������<��e\���6���'�ѥG�v���>k�-��mi������#$b^`F޹��ݾ`��eQh��N�]Ec|��v�ɻ�X�Ո���X�-(L�\��^�눤�`0X�-Lx/\;%�|v/�Y�wi�6�brg=�|=1wt�ȹ��}��Z��'oQ��p��5��X� ��S�|.��S67npi�9=�X������2�o�v5�k��f�
�u�	H�f�я[q~�%�1�|�x�}.|F,�{�]��'h֕(�6T��1��Q�H��ʚo��}��wF��S)ӛ�-�,�K~���Q	�V����58qa݉��^āĺ84��>��e'ǜ���7@�L'�ճeM�6�"~�Қ������c%G�����<�� SY;�3l��k��n��x�v�:�y��}������	#���8v��Aȁl�\^���k@C8O�W��iP�c8?ס��ͬ�����3�8�1�N�(,�����#@%�g�����_ƅ���@��W�� n�l"r)�wW���/ע{��!*�
̋)��5�F��f�ݢ�1��!V˷��V�r&��Fg/K��ӄ�����ʾ��n�J�Z|S�]ЇȆ�*��Vۄj���X�qؤ}\�/��%�4`2�}��l�h�����������'�ePD�V.�׿n)<�Ϻ饐٩Lw���b�r�~_@vϻ'��)M�+m���Y"���k���-L�q�O݋ɬ�"}r�ja�C����q2�(���r�}��[I|�ٺu���ka��_�|�^���sXwH^;/Q���I�Z��+�M����R����ʁ딻�`�c�5��cyA�Ϸ9{��-�6P/���M�	��|��{Q�Uec��Jyo~�f���r��z�W�T��tUgcx3� ��do�_���g�WQR�R;�Ď}��hK�t�7̑ٽ��j��j�K4��=��;��q8�,&�j=��c��v��5�⸭�U9N�m�P��XE��5�z���F7|Ŝc,�i!ox25��&]f����]܋p���j�	E{�h3*j��w˕#�2�g���u����v!����2��.�g�,q��E,/�4�<�ݙ�IjX�t����������l!���E�jyU���� ̮wlKq�Fs4��h�v���h�b����8�Z�E:�r���a��Q�zʲ�-3��f�Xocz����jr:(���_+s�c��!X��'k�z2e��f�fB��+��c��+��ˮ����/�ϩC�tě�af�cF��� [G�����dI!엯�k-�x���S��z�'��g-�Y��Ftb ��R�t�j��"�=b�e��ሢ�
��Y+���~^L�j�%g*Ūz VB@8�qۆ3�/�Xu�}Z�.����X�kXv��>���z��G�{l�ҁ7�q��g�ׅ=�6k�,&�\՝y�QXa���a�B�Muɽǲ��K�N��v�q�̘�����/*�*姤��KKr�2���- 
B�3��ݿ�kt�����/]���X�r7W],��Tmwb�Z�~�7��'x����c��R��\�E%�L[힅��T������>Rv�t�[1���5'{��?թ%�ic N�o�V�F���Bl���;��У������"С���}�\
��xMM4�%/��|��:��fKeqX��D_k��� 5����p)�1RD�3�_��A��j�պ`�_�5.=ZYY�xW=�p���~���n���E�sW�s�C�Z^���-?X�uv���|k'#����gn�8�7�MC-I{vi�]�iA��s%ļ��(ev~�Fނn�d������Qg�?!�ķ~s?���z��ֆ�P�9���S�?[��E�12��)U�]#�n}/�vCN���U�֗�
�;֭o/?�^o���3n�q�@r��,��5�0�ʭU	�
�`����%�rn��x�b���uE�Ȭ|%V���}�p���O���a�z�j�W����m�
�g��e�%����Ke3��5��yĚ��Aq��؃/%�-�_o�^cg�g`}m���0շ��>6�R!����2�K(���ĭ�*P����`pZѐ2���������j%��(�47Ìhz��!����I�gw���V�k��(H=p�q���?�KXv�:�a}�=�T|��>4R�9as��&A+���{�݆�^��aj�U����*j�xWN|/���B^*��� u.T�q,��<������@J�p�T;Ȗ�����=vZ%|�_d�t<lZ+y4#���7����SO�
^s?3.g�jRs'Z�C��B#�����^4	Q?�=5Qn�;�UP��q:�+Ui˔[�g�W"��̘?��<Ş��Z�i���|���2��r9ǜ��Ŕlz8������6*��L�1��bA�В���5q��ֆ��݇FL�~��L�`���_�1�F?��7?����'~]˖a�7��7�b�0����c�>�;�J��i�Gf���-�t��q�ϭ�Ľp�~��}�n/$N?�V�;׷��, j�C9��UO���=f��,ٮ��i�����¹�Ae���T�G-GН�L���Re�(HK��2��X]}�p�wf�-Z� ���N�T߄��#/���/�g�eK�˫��71i�ƣ,�"�� s���#��=7�/���[�j��BO����f�+ӳ�k��*n/x9������떺����uDTdF�����F��ә1WU>O3���	k�_oh��/CZ�z�%����Tţ���_�E��n�t�� ޜ�P���"�!3hb��"C�w�����sF�1@�K�W�L��kݽq�N/�b ����/�C��s���nCi��_��δ`W׎�&Ep�p��k걹3���۲�z�>�R�����i��g:d)U+�i�a�.v��H#��l�'Z���B�+����pf��&�/]���z��O .��
Ep�c��$"J���b����P�֣J���}��w}��(�M��`��{pa�Ũ 5k����9�n H$�kL,ɸ'�����S�����aViN�w��*��@��SxWz���^3���4,08:�踌������꥘��H��������!�a8
��ouK�e>�(X�:�w��=��V��= G�K����'}od��6m��8�;�b�E�� �-�4f�̜t�|Y�4KQ�cG��v��6r�Rv�Ӡ�ԮQ=� o3�й�@�@*$���߂(<aN �_��Ш�#?���w��|cj�w��M/��H��j�G�j��0��~��!8�����4n'[U,��^�R�%h�PwYK^>�`(�������T:M~�n���;��b�`��8�h��*�=�ꀾ�f��Er"���X�x��6���3B�/�%��~<�)�a$\��/���M�;�a�֗�ɣd��Z�m�5����8�\��SK<��	ELT����=dk�T�u�̣E~��% ��(
�%���py*��Vj��h��r�G�r�Vb=��qo�k�ޑ��s'r�����gy_Ќj��[������9�-��D˷CZݍ͈��Ħ��o��ͦ�操�b�����ćb� 8��I_A�F�� � Q�O�l�r`7s��i�ڳژ�,U�7�Y�_�r��d��<�:v�P�.���l�Z�O\� ��9h�Fm�异���V&Krm���ȷ�Y�! b����47�K1l4h�2�3�Ȟ��.^�V5+ˀ*�k�� x�eb��D�<ܰS�;f����ݫuЕ��~��ӗ2�k�5}ƊR��f�~�����`���h��|�H�'��!9A���X�x"�5�	���`U�c<�xԷ�V^v:��栬�L����-NX/n��#�UϬ�bu�d���@���ݎ�[qep&�Ku�S)üb�����P5<���L���as��M������'���U��3ŏG2��7AW("����ٯK��ag�b�u�|�X�A����nb"gg�1u�!�DIݑ4%�!��f���Q��T��Wv(��d����N��b��U{�X�L���G��{��'��!���&���QMt�h+j��f�٪/����QXK�=�Ė���Ȉ���U�3�<m��⿗�+����M�WU!ۍ[�
�ys%j���o�%3�X�����o���~%��h?SX[!�(�s�Ķȣ�F�m���-�*�޻�+r ʀ�T���cΜ���D�R'|C/q
��t2p�v�<��6� �����J�v��f���;#15��.�Ӑw�Z��(��I^D���r���N���Ҥ����=��C�����Ư�%c��1����C�r�cS�(��D˭�_�
�\�G���v�h%������ �/��7
@�7x�S�@ׅg�}z�?��Q��D��]z�Ђ������!���?{r�,s�^��1E����7@]�o:.�Qn&cY���Dr{�Ù.\jIU���/EX��y�|����3�+�/�Gf�,����nڵ,��qf �ׂKu�*��{o3�����O��{O�����zq��\.V�?����k��ꬪF�{j�.`?f�*M%^��u[p�4�U������	���a�LJ�m�B��;X�9ǰjC/�*P'A���S��X=]w���~|X\��a5�o���BӸ��7�e�nUN��LY_B��_J^���j��S�F�g�錃A��k��*g�d�SS�g�,*���?�����>-�����AZX��D����%G�O!Lɛ�A�Ѷn�z�����*XI�V�E���;���T��K�V�%!P�e�g\��s�/�����GV��+����Ԕ�\?D�$�B��nn���'/��U���ȩs�����V(�?�����H��
بӱ6�P���Y�6���#7���bP�{K�ҏ��6�i�Bm� 
�Vo)ON�7��� ��� ���(�L)H�U/�^��Q
AO�iW�Y�'K01I�&��O��^��3��;���G���Ws\�Q����40�0�-;7]\��!ʹ��5j���;���vZY"��.o��9/j��NEE6j�����OM��Ÿ��Q���t�N�A��Sa�0�z�c׊Y2?N��8�x	����?V�31:r'G���	��3l�� "��F�D��&>r��W����Q��mT��W�G2��§v',튚�nKڽ)n_ pR�m�gc��n5hw�T��xiR1'�B����r�<�ov��MOl���~CϚ�<A���H�����5�g��3���f�q5_#�F�Uj�p�{VIB��8��"p{?!9�+���f���v�>`�s��R�@�[N����3d���/jӖ���I/��fs^^e㒁8_����<Մ�6� 8�HH����_v�!�*DP�/�|�r~L\}|����2գ�+�ჩ�9��TV^�f`�q���l'R��?[j<:�ʄ�
G��î��0��jS>\����O��T5붕��gC���oӟQ"1�n9���"�VX��ɇ�0x�`��4y5���������ˢ�k^� [��l��~�/p�S���-+���7\�|?r�V-��;9��[Y	�{7"�1�ׅZ;wy��!�KK�{p:������(���ؾA%��iI���¹�M���|�p�E�ؑE��3�K�U^AL�c���b��1G��_f�Gh�a�ߜ��'L/����FT-O�o����4:�"f,�v5�eL_�w�9X�Z'�y�Xz�nk�86��w��N�-?�g$&`̃��U�WcOJA�kR��7d�'X�Y�at����:�Ծkp���bc)w��v�e�S�PC�Nm�*atdf�N4�k�m; ��<H��@�����/j�0 �_�U��LW<� al+<��b�q~f�bmNL[��)<��[V�޿����m��}�J�\Ȗ��)���nY���`q����֙d������pnAǔu|��@k�8���W
S��7y
l�F�qE��F�sA6)9]���6�F���W��K;,�U :ǖ]�{��+�?�+�HG,��W�����ۥ?ױ<n��i�
��[ݵ�gJ�����Ѳ�0l��R����n�?����Tޣ���K�PU�5ʚH��l܅�k�\�mTyRՈ���@�J�fml9����Ed.� ����Q���uX4������魣 �mnU���w��Vn��~�c.=�:�-[�ܐ`br�{	C���Е�=�K��@��*��mT��j��y>M2�J��I�s\/>R�����]-k 6|--�&`_��u�U�5��ʽE�S�ק��m�ODn����R� 򾧫[�Kq;�i[+��R���~�&�]�zؓvC֙��!h�>�\!L�Ղ��w5+R��t�O�C���m��s�����'�W���ʭ�8��s'kpӈI=��A�+��o� ��AN�[�As�Yؕ0ְj���D����i����?�Ҏ��I�7]�1s�P�e��4�����b�˵qԇA �+��������Y�q)d2�It�{[X�9���c5%������1"�=q�݊�{���*��K��W8���:y�y�.�x�H�����{;��>1ͨ��0�9�W����E<Qp����{IK�jJZ�Ӓǯ�-��=z��):j�}M捜ͥc����IE +}0�J\uPҒ��u;}�D '���3��G'���k��3��>�e��,��䱡�9r���(��(Hi@0�*���, �ѱ/t��=�iN���ɅY�f�𷑤�w����ӍY�zB?Os��nM�%���'!�L��	��lJ���耰�O�d�m�qy���t�'	A���آ����	�z2���e�l����d��֏��^+�{#)���7����:�L֧�۠JzÏj���i��q�L�R�q'njDD�ce�z��ԏ�{j��*ukwK �g�S܍4����V��c9�[�X�I�(99 s��������ӳ˥0�K�?�����/,�_� �g��вi�M8^�-7~������KHI�ȝn�v�P^i::�9���Pә![�_h,��B��7��زU�9���vsK�f�=)T0��zl/ݤʪ�R[`�����h���b�&�p593<I�>#�n�bC=^��B5��3��`�����R����L�}C��4��� M��_�_�{c����2\:w(=L� :�ĔQ������ی�7Ъ�/PU�1�����] ���,�U%bF��Zl���㳲�x<��� ��|�����ڋ:Ú�_���"tk6/'R���PU)_��g��8%eOY�����������ˣ�+��������?|z���'�F2��H0 ٕ�S��øv�D�5��HH�;�xrȧ�	�K ƞ�L����[hM\2BQyT�Y�c�3��6�H'v;*�g�	f�"�3&�	�mtٿDN�.��~u�qpf����;cƶОS.p�E���K�=��8~�;��n9������`��ɦ�u��:u�7c���{son3ވGJ0}�0uz�����KGOi�Mj����4s�K'�2��oʩ�Lb���4)'��"a�L�K*m�*'�tE^�-�]��_ߦ����jJ��c�����}�^� �Q��NEA@����* --6�G
H#0F�4��5���������9��}]��;��r65u�t���W�@84��`�,�`!j�������u ����ɪF���O��&X�Z�{��r�3�8�_�6��R�nY�0ft|����6{E7��� Hn�9��:r���˒�ht�����A�( gS������1�;���������#.��O�؅!)IH�y��:�2׈Yg�]�
l�8ÿ��B�K�jZ~��)�GT�ӡ܂%+R6��9�Ivܓ-���S�����>�f��]��#�>������$a��MiN$�k?��(�e.4U��9�ǝ+�]��ҹ��6'�r���[w��2/bAp��f��|�����x��A�@��5��x!���Уd�dT����� U��A�E�$c�^��-ω*_���p���f�b;d4���θ����t��\��?�½���`(�A9R�oK\�	��%��Tx<�4��\��Y����}�Xc�6����!��W��:���g_®�"���<N-z:E�{�0o�q����d��l�y���rVSܩ���BWח�	�{��ǯKfe�0�7�o�*�o�����R�V�]L�6<s�ˀ�ΰ��"���(�@q��_�r5\��}6�Uk�Q�?�f� �a<>��i_�@�@�<��[��m���,L�Ll�A~���O����\#��W�o���J�cm�˾��?_d�a�+�oQ���Qb�{��%!xx�e�;������f�pm/e_�_y�U5�gD�"^�\�堉̨���=���RD-�8�R��m��>ŕB��9:��"Yv��%ڼI׋��ع��:����|�(X�a:��sVJò��s�t��"���8�s�LSV���f& #�:�L��-�ʏ"Q�PRV�A�/���� �/0)�u�X�u��%�rce�ga�8nPG��:��y&��� #�<&r��&�f�{�b"9�4��	��ߒI@�ʚ�j�:'L�]�a7�	��}ԟ��RT?�㯍��T�&�rԢh�������zsmO6"=0�J"���"��ASz:6K�v�І�oܓ��;7K�R/ђ��Db�������>�}[�C��wPz/����ݒ����ۋ,�Z�W�r� �	h���Z_��.�l���Q�K~q26%�k�c��z5���ҲGu�M���;�fi�4._��l���
�Xl�A`��8� ��c�/:�(!�OF��*���ǘ|�H��$_R+�	��n4���*$d�w��ϛ����F�}��2��$����!�a;5۽�R������>r�n�Q$����������S=v��[��Re".c�B�JR9�h��F#��I_������ʩ�7~���ҋ��`���(URVN�[��ܺ�Q��TJ���Mn���i�40����9�Qr{ͩ�Umڝ��qL.r����Ԇ���w������X~�2��AkBl���>!]6*�<]D@*39�X�k�!q�!�8��2�������b�b��fjm<�V_/��/�)�S�Ȥ���Gz@���T�ޟ)�\UzU��p���_�`���Jc�s��5��MbFM���RZT�$���n|I����&k�N�̦�x����:HMzњ��g������B����㺵��*L}��Ě-��+7
�ءӥ�]-k<7
����JC#u�eҭՌ"S�e�<�����K���Ͷf�="��l~�Ĵ�ӳ�?9hSI��uY_a��QC��c�1l�8%�Ùђ��mC�Ò_�^�f���%JaU���|kyZV��>P�K'y�-~
���B����¬i@���|�s���\UBK*�0�F�}��������u0,Z�*Q���N^���1��N�.ZkR[�u���L_��_�_Wt��5}tƐ�[���C1]yT�HŨ�r���u͍�0��]�k��:��c
m�������%�x��=�IU�8N�B:|�@S�x��wF V-��%w��#�p����3�^���y�WT$��#��06݉o�Ei"O��*�R�3�9|��j��lo��[p�����ʟ9o���]V�&k%�^�HY?5��&���ؠxt6O�?-��:�S��Ǵ�8@���W*l ��w�5�IKd�-�q�(��-p��jw�vI2`�َK>�D�!A�II��;b�7���_j
�UZ�a���7����)��4ɭm�Vٗ٩��y6�7l�(谞�§B|��Q�Y!S�H7*O��:8$�!��7�ڟ���U����D�o���}�,ub-�k�'�oh��:��8�І z4����<���j�q�Ya�ٯ��%|hD��c��鯎+wӬ�P��T�D'
zC�K���~�m�Ճi�����X��빜
���SCi�� `�@�i

0�o�åڮ�V�I�ORLO%[��Zhk�)�l&�:|�yRº8Mݖ�(IF���}V���e�M��'�����Q�`.e��z�r��W���JyNg�kE�7x-�h	���G����}�X,�=:{T3X�)=5�}��'oӘ�X�&n;o�E�7(�J��x'�[�� ?�������D0r�?������F��|E��EC��];¥~��>Ɏg�pz�`U �׮�s�z"gm;�6���C���U�$�5��{<.��r���|y��(V�z��_�	{������fvX���A �[�$]9����y�
�J�g����?�>�=���^��W�&U���?cA���e����M��7u��.���U޵�j��kT62���]�el�nNl�MMK��^OD>^2����<��uz7(@�Җ�$�E��[\�`4��sƩI{{.ߞ�	+�,=j�p?���<o����|X�}���?���@\��􎷣ZD�o��7�"mi�Yd\��R��G�A�����v\���gUnv�և��t#��i DC��61e�<F]��8O�S�>z�s.e]�|�[O�p�͝�<�ӂ��$]$鑈�J-�����3eBȞ��<ChA&�-�3��9�_��1�Sc	_D�i�jW-;!a\�R�!\��6�r��6�R��u�^J����'>e$u��k�>RP[T�j�R'X�-���K����a�����}��"	�������e��uD��,ye�������F��V�m�Y�8ឤ������6�փX��i��b��f��iW��T�fr���N����P���# �������8ں3.^Ќf��N��K��I��2�vV�--i5�z*G��K��nO��JJfS�TZ��i�F-&	j�����Y�"�ѫ�t9�;�(�b�>��@n������b�%�~7�����s ������k�"��a�Kz��V�l�_�p,��w�V6&�� ԓ�M+�t�yvD��H����*��$3���z�/VP��4��M5*�!X��n�12��7���j!ۯhz��*�v�\�������g���
��e'yPv��3��q����Us��;1?��k����W��>@e���:y��а����5��/\9�f�A�jɏ:���OU����N7KL2������E,�QX<Qw]݇��/������4'�G��eO�S<򢞤�4xIVi��Gv�_T�N�/��<�p�3�GI����j7�NN�U�ND���t��yq��צĪ���ZC��9Y�ւCS��"�[����?�iR�A�5����Ü�:���L��c�C����gl���|�.��ζ81�)P�yu��T9(>߬�����1����7$�N�s����?����s���=��|������g��N5�" �I�7��	�7���8oZ�g�j�ǝ�&�R�T�l�i܍�w�g����!�y�n6�u�$Į�9�I
{��{y�#��h�5��#�U�Q�L���?��*�����uw�����`*����yW���T��5m<Q�����/��a���ݵj����w<J#w��hev`�r�D�� a�|���>� ��r��aT�|����.΂�췩��e�5
���!���:��b�쳝"P�v����T��aU���"���Z�+Dk	7���_�I�8�D����3ix�%����V+�!���σ|�C����K�:^�;j `�:���a�7�w�B���.��>yD�60N���F�?��w���5J'�������jS�̃5َO�3���]߿2���ǖ�+l�Q�s�;��:@>��h�B�}V�\������k�SK�ӧ���n�ɦ+o��W�Ig����]�\U�7����b�>m0?l����7�U�L���&�����9��`mk±�w��'2^�i��n��d�����Nw6����6�E(�-B��$�})��
���]�n���}'���o�>>��E�-�(�p/=D������¿��ƕ��
����+I`�AS����zvKa�/0-���~\�\1��xߢ��'�T!���29_����NJ�ޮ�f�Oڧ�=��H�Z����)���O��=
�F�1�$�d�X5ͷ�o-h�����8�1���}�.����KC���~3:���:賂��%�z���3����2.P_�ܡ �e�؛�1^K�K��Z����c"�C�E[uY�	ț@'F`!EE`6�vRU�����N:�u�����ƙ������1Š_��|u��H�QMM�T�z�k�L�W���J��6C����Ǳ�2I��d�,"����~���g�T��#N�`����?�Wԇ�`���	O�����ģ溛�ϑ��Z�}2��g��~��m�&e2���;;v�%=S7�+ۺf���5�F��-���	L��l�v�ëm2�&���a�r4ɶ�������n_b:��H�y1�BH�L\�����L��#>��1_+M����[�>��x�����V�^��];⧨�J�'f��2�=1
3�\��d�U�σH�K� tя�`::�}�K��榈+^l]1o�2�-��G���g_`���4��Q����x�����b��}T��!W�yò*r��[�u��&�2åoa�{9ԋ1 C���pST�M���س��+*������q�.�wĽ�[���Vc�?��|)�5֗Q&l�_��H,���☪TdW���鳲�����0��>����5�$|jr�ͼ��Ds��)���G~��f����җi|�����|8�$6?l�A�┛E��Qs�� ���0%1G��s��D��>QT�O�#�y\�N���v�"�ꓚ�O&zCL����w��j�a����ԯV4��U��D�u
 ��u�)�x,�7�n�X׭d��3M����6�����BY�}�\��qu3��&�("Թ��3��L�0m��V�!��T��x��8�?�]�a�oV>�u�+$f�̗���89�(O`�¹���ײ�riD���󇫤��>����@#e��z(��L��q���g�B���e|+����QQw!���C��~[_�=��:8���KqEq����'uc�Z���..��c�$6�M��ٽhބ��.�@�j�y���s�A=�@�g�
�>Q�@�:��'U�)q��:c0�L����mTv��;%��5�ݎ��-�k,�YKIY�^�eJ|E�9W4
&b���I+�;xӶ��.�w�x�m�/��5t��H���aI��P�y�HPA�wV]��+͡<,$�!�k�n���8���"��q����4�dwm'���c�T�W�~&a9�KۚU�tVE�J�=�y:���1r�%����f�XėI�'�#��w�P������~��_�Wˬ��$Ɖ�9���|�Y����T�|�V�B�H��jL�I�:���2FKTfK���g�@w2������=��F^�L~I��C��l�K�����#�B>�C�h5A�-RTa]��3�����ⲣve
��98�v�U42�韗D}��%o�x(���+���.�ĕ+�}V�F��I��7}H0�	D�mf^u�7�$jC^�J�|dk����,L>l
�\i[�����]0.|ӁY�I)u)�&�C�7*6kf��K ���s�9�m�s�͢��}��K�<_��$��*� �`��7�nkoW��濼Z�_���oӓ�jDUX�����* _(K�l߸V�n!��9���z>8�O�ͨsw�N]��U�Cm�C�����A3�]��x� I�_4gF���ݙ���*\��ی[Ww�A��	��ˡ��9_�KD�����&�}Fu�1�_/a��Ru|l,%��%������_�=�n�c�{w�6`{�7�7,�n�n�k�&Jg��V���ZM���O9#�0��M�ʿ�Ĵ���� R���T�����)?�ؙ-P��g�3�� ?��o�ݥ�G!���ϰ�3	��O����۟ʋ��&М���wb�&����+��V�D�$Z賳��]n��SdX��Μ�
�GѬ�[���S�F��1�J;�"���3p��ﮐff[��͍��#n~�M�k�̈́��)�3�m���He��R�ؿv�	+�Wz�a�]��o��ƶ�����5Mh�`�h��x�3Q@�$�,��[���;�:�K�<��#4�����%uѫ�t��4���B}�܋�a�+�\!`�C.�݉�ڕ�,��N��x�-W�-���o:ˀ�"�jZV|��2)����X��Q�������'X�'�A�t.���b�K`3��o<�lnM/Q�Z�͎o�+�$�h�S�7�5K�(.��!���X��q0	��|!��2Ð�l����:Y�J����>~+���ٝ��}q���!���� /3o�pR�m��k8߻$>_ej� �Xl�]2{I7� �\��9���CPJ���=)�v3�	��ԉ�~�:���@�h3�Yȫ�>�^�_�I 䙃U���z2�T�����H�1d (��8Og�11�M�����[��7 _�FF����p7�רQ���p3����Eyԍ�4eM�����^I�/���m�Q�N�Ö��t�s�]T���C�;������4ű�\Kpx�O�Wʢ���a���dQ8BG�#�~Q�9��E��Cթ鲱ޜ�O���U���vl��L�A6�7d6�~��^�'�A$�ƝVY^81&m8x�N��\{&B���>����7G����5��v[���*�M���qㆅ~ܯ <����TC��z��4�^;$��q��iԎO[���?ɬL���0[�
&��/�G�vv����z��a�y�S�DeG��DW���)�����9K�x�t��T��UX��l��
�A{/�յ���t$�"������>=���?�{
��o�υ&���..���x��3�m��i�(����ꜜa���2�}�dR+���(Ĉ�SR��,��K���*E,%�S�ɫ`��nfN0�;y��l_���
��S�7�;RB��Q��BZ����ڂ�DQ2a��^���Jr-�;V���c�ݖ~��E~<���PL/��(��=��k�T�<>ؐ�����(^m����b)��D��TN�M%��g����`{$-MR�ݻ�GC#ȃJ�Y:`��!�D}Q�\�;؈^;l�mR��[s����:�mu�C�ۺ�e-GGX	�F�����2*��#��d�~= ��Hxm��N���!���	Ĺ�9�V��V2frziGWzl�D���=�I�����:뽕ʵ6w(*LYw�ag���<������ņ�t��rרּ����ݱ�C���`
*Bۀda�?D�;׉\μV�A�PJ��'%Sd\i7vo����	kDS���X������x��3��qƖ��ǣ^H�(�e����ӟ�����W~7X�?�5<��gj��޴��M��3�4��]�T�Za��r���P��f�x_x��9_�Xh8���\�ϴľ�~����_��K�	a�|l�_\^x������e���V�	����俕�Ư�S�)5��9<9[w�o��m��B�v����S��{9�|�?���}��H��m�+��W.�֞R�r�&�z> `'�u�p&2P��&%���+i����@#'*7�#|]\J����%1y���UB�&�TI���s<�]ȡ�x�c/��m�����֍�@�ԣ�O��s���/27�����f�#R�e��=W�η�4��7e��M�a��/ۦ�Qz3�o����'��z��mMS��-�܃�wD��̓���+E�!�ƫ��t͜C��r��oNTu�khDrrHI�.���hd���8�rv��dA�?�����}�y�uǧ-�EY�[��8�l�����am^���G���+�(DxhD��O��,���ޤ��y����"��v-t��r��*�>�v�U�;��n�C�r?�m��7)I)ޗ��2�7䍱����(��wԟ�~N�y�U�#�͋����K����"kY��z�a��!2U8B�B����?B�^4}��ă�^Z,�<[��:W�'���H��YՌ؁�V��ߕ���v�Uvƺ��
2��PD�^L�}�jtqZ�T@
�����Z����ʨ�5b��}���~[�$܂-�Mtϫ��`^��Bx`�=9'��O�'e4a�9���"  ���Oq�vil����/]��|U_�Ѐ)��Ѩ���DQ��r�f���:��Ŝ�F���[7��ۘ�+Jy���m�_�f:�����N��1���/��'�R��v�v����`����A�oޟ�ڡ(�	R����q��zfB���¶�,��M_�G�)�V�/ㄽR�t3����s�iڦ���;g�����҄�M��p�7�����L��}�Yo�p �OH�q�M@*٤כDғg�¹���}��O[؈/�+�ׯ1A�G	r�"c1���m1��ʟ��R�J=^�+9��װ���}�fj09G'�QO����kd���`���tȣ	H��uD׸��D�;;5D�	I=�U+�uޥ�o�d�z���4y��/��d瑭#�q�j�Q}0�~`2$N�Y�Ii,�ֱ�dԹ���'��##�%}���d�[߃�'�Jis;�m�K��?2C���R�d?k���W�v�EZl�Ȋ$��=|�4��H��\�H~�\�;�FA*�C������\(}��$�6us3&&�b�S�o�<�3_e���$�#�����ա����L�(�I�$�s;�ո���_����ә���
����k��1D|�T%��bٸ��ިq������h�F�q²�Ҵ_
t0{F�rҬ���BK��#���,��Ù��!^@e��j���l�FW������*��g���=���:�sY@���S�)~Ŏؽ|K��4����[B�W�CZ+�����K�����/�6�/��T�����c�s UWuP�^��B �����M��T8Dt�P� �H��&��\��us��RZ�2l�L��Iy�[�~����DЀ0*���G+>�L3rv���H�8l'�����=�Ө�(���L�Hظ� !�V��3o�)���X������-.RUx�E���杞�e��S��"3;�����0�B{�"t���|qy�[�}Ǥ��:�S}�N�Nw���!*JV ��ڍ$rXO�|�w*�d9������ǃ�>�댿m���[	��.L�\tx��aO4���b�Ґ�'���1�<���ࣼL�:����orI����DK�9H�1�Lί������k��Y����ua�M�������8��v��i�BB��;B�%ލ�b+ˣ�o�r�}�e>0∎��5u�)��g�+YoG����1N���:fB��!�{0	r�〢�;|#�|#[W��(�ܽH��6��@��). ����&&��K�����+�z����'��yQj��@�GRۢ;Y��-yXE����B�j��D�Xk^8m���I,5P�Ra����0��g��m�͏V2�>u�ʣ+�/��f��}[�3�L;�"Y�6���U����
j�Hy���p�d�&qV-&j^u[�ie�v���iD �ʴd�v;���'�0�&l�:W��\b�G��D�j�H�kX�E�l�f�V�2Sݲބ��l���v��GA/gh6ꢫ�3���e��â���آ��-����G�'�ag����)߸�g���5�ˏw&N�wI�>#?[舚�A��3D�/�­?x`��Ӗ�:1p!�g�j��ک���r%/3f�Ԍ��z�_F�d���@��$����E�X9x6���%&4s�`ֵ���:�L��.9Y�a<�N)x/�*l��Ku�����>����ŭMb����{l%�]� I�ܿ*9Ձ�&��_�t�IL2�5��#��e��yQC�Z���fG����䮼����2���Í���B�~���? ����A��%6%�QS ��c�|��2�K5��s:S��&�}RM:Rz|�zt��.Y��]�,�mv�Gei�'V�;kh����x�Kx.�\�Q��<&k��ɫ3���Y*��n�U�x�`i�K�zl5�}���ڭm����s������v�gl�sŶ�i�V��������B)��Z�PEw7�h�s��?�5�����kq�8���b�ʁ�w�Pw�"W�� �I�����i	�)�6^�k��=��u�Z���I�A����0U&&=�q�B��E�C�,佽K�Ͳ�(�14Bc�-F��G[<'��~�.�N�rre�>g^��KG�� �Cb[�;�P6_�z��A.��۴�х�deƇI�"�2Bʏ�{��e�L�魷b�տ�B�J���z�8c}ٳv���3Ӷv�u�q¶�@�|��֝�����e�IJ�Ju R���E��n��C�m�צ�������ȕ�VD�t�&c���.���g��z�"�S��Ls��ΕUt( "��u��7�ѐP�p (.� �J�UJK:!�o �~�1��_=3���=0��X���qNHB.k�G
J��=�Pc� $0����|3ǽ-.�먜&�T�FU� 1��zii
P���5Y���I��S$ʰ2��`�U�o�� üH���;�@R{��_ȴP�iv�L5+��F���sY{�93�L�������V#��ή�E��l�Oh ��N���Q�t<k��W�ܣ�h
��ARD���G��������qʶ��[���\ӂ�o`�~��|�����PG,vm�G�Z�t�k�2�lK|y2�7��ɝ���Շ�����?����:dgq�W52�pJ�q
Kg������+�����\>�`�����s��&����"�c�,S�G���?�H{�۟u�i�5jj~��;�M�w�t,���6pL�ߨ��94�O�|��}��)jW9yp��G|���kv���}�8c�>�F��7ũ�(�Cqm{���7r+@%�&�G<?�&�*]�"/O�> j���Q�޴�@8�/��Q�6���x�0LMI�N1��3<w��I�@��5^��i��вno7�M���s�{����	>��t_#م��Ks���.6��M}�*2�K���i��%ғ�	w�=��,�(�Z�ܵ_�H�k95~�� ,2��9����^J��b�3.�Rr��P�OmO�:$F�G�T�'�x,j|򥡫�h�p Y�	<(+��0b���+�B��BPU�.b ���`��fX�.�@C����+����}u��2R��)�M<?��CP��m����H��ba�jЄ�7��+��U@���L��Y�����4�>=)
�۝{���È�� ��J s*+G���0�z��ǲt�EOYۄ|5�,�9��'����,X
��\���=C���˽)�Rԣ��"����(63�Jk��V�s_�����V��{����ks]��2���v)��]}��FH&�:!Ȁ].��s҅�yp�1S�ֺO�BQ|����%j��Mȧt̸OOd������e{���8�3aǁ|���d̪�GH)�T=���I�K&y��j����2���E�x���~�QĮ�|��1Mo�jՌ�����&�[�u_��G���l�!�w�0 �h�c��j��_���ؗ9LF� bp#C�M.�ъ��|��U��N��i?�05�� D@���(N�I��ȉ��o�\OW�^ե��2�6���)$�LoJo�����-uD4��+�l�+���!�#��'pFӴV��e�1etӤ�I�������RMj�t�/��$*!���>4Ea%�[k#z�#�n��o)�X���
�@�n�;R_�ḻJ�3^&u�Þ���������z��)�h�"��}B����ep�2���~��\���"��`�������m�s[�)qJ�@3w�6�C����#�ϽZ�+�},�U�ֽ����**���k.���G�ۓ�lc#��93��+/ݍ�Q}��!��.�skQ!D��V�)9Q�Q&����8OL��c�2���b�~|�:<��Y-..�� s*@![O��+�*�����D��"S�}�^v�eQ��P��PW��C���I��j^ȭk���9�+�ۚk;ĳ����+m�������������>!�|F��O*0�g)P���+����}' I> �C��z΍���w�߷B�:�-,�9������m��y�F6~K$��q���ٽ�S^*�Y6^��~>h���^Y�to��I��ndG����\�V���q�*Sg�����ׯ>��(r����}x\ϳd"�Y;v1�=���l��9[ԋ;�S|ο�r���IJ�7S������G���06��[	����x���BS䀺ӜrU� p(e���ґS��A��D���/�2_>Pؔ�*�h��`�� S�l��C�A&,�܊�
���6�h9����w
*9�L�tz���D��4�r�I�Q��K��2���f��R��,I`�D�UVY}��|`��N�7��V֎?�`\�zdT�CWl�=ބ|��/Lk3���s<��O`Y�|������J�<[_�D�+��w��"�>��N�ℚ��v���T�{��P��5!�>v��S,�4�w�݋ 1х�&"�#��Wۗ���]Xd���L���C�9�Ӑ����]������A����,4*f)(���l^^P{��h�`j�A�̦��w����
n�5���D'�Sgw�ؑE���%���;@8n�`rf�z�ܬL�;�Ɲsք�$X�W�+�H>�xp:��9�]����}���%�%4mB����Gn:��/!S��FNjA�תz�$N^)`N�Y4���<Ӛ:]B�'��a��AJ4+J:P�[�s/^�?H0y��lB�v��?��vP�T��� ��/+qii�w�VTTP��~�������1D��k�׺�Fְ10�v�>\��Rl�ISg�X���p~r�-`����QT��Q��R����7-�$|���^�h
�q�}�[�[@m0O�^�-��T�F���C&x���Ip�j�L_Z���k���A�q}�x� �?�����{���-4ҽ�����-E��ĕ)����m�<��Guz\'�9	�+�u��J`�SYG��;��S��v�ҿ��oR5���2�TMk��:����S�8�&�+n�09N�O'�����4�kƯ��$ӛB2�5Vr#�1��<�(��Vt�|BYM��&��\ƶ+ޥ��Vu��H��Q�!aj(s�E���Ǚ
|'˙� o@HH�Q��s"m/�aX\��"��y_�Ae����w�(t��;��]IAȇQ4I�l��	���|p3ӯ�����q�3��B�s��Q!|T"��ZC��w)7.}��&���I}y����V�����D}�?����k~�.eϹ��Y���9f�7D��OCnR[V^BD"P�ޓ��|��D��^���h�?s(N(I���&��H6�q�{�|�n{S�ZP`�?�
��%�1� >߆Jy�"c�K�tO$/R�_�g6�u�V�c[>��4�i؆�7<�qsu��?�PXÏ�yō��㻖���=�ma�A~�=��=�1����b�%m����xU�ϵ�f��%��^S.��Ɍ���0憈7�5�g�a"1z5��dqm�kw[-��jkk����[1�x��3lG�m�wH��(91���S�C��Ƚ`$�Y�T������/��i��T��-M��%�bb��	C�� ��f�7�7 v�㺆��H�*鰎����)u�����e��D���*�`�����37��Q6��Z������rﲖ"����1(��v�c��*n��?��
!���`�W@�����3�q,t5��m@��8N�����nn���P���	0�=q␯S쇿���Q����rZ/Xds���(DT�:G�8�����S�Ȉ�ټ�7ēm�S�|�y���7u��i-y�1N��7��͌�BH�>��mj`.R�-x�ˬ�=���f�ws�q�����U���T���W���(� �abj��dr��1Q��V¢Ϯ@��E�UA"�b|�B;*EǱ�U�H ��@�"����ʺ7�M	{q������*%�8	������I�m`5 8��~���ؽ�RW���[���e�:���qG8h��G�eQI���Ô���_dֵ��e�*�g�~�����b�+V2�R��=.���©!����̐:��m{N�.4�Rxg�z�'��t�J���8�z̢�m:�H��8�L���t2�ǼEhro�0� u3�k�Mr�K �ux^^���B|��J��|�4�?-�D��c/���t+�6�)VZ�񯚞1{7y��?�{Lс��̿��RN�A�6�?͚�F�e����a�T���e$�8��l	1��a���՘�de��i����r����ͦ����t&�Ef��<���Q(��5a1~�[3�Ȇ���e[k���wU 2�����d���:��יD����.��[I�7>���h�`|�8�#$����V���F��櫘Y�hu/D0Շ�#��%��oQ��A�}�{������i��8�ؔ��2V2b����v<�}�>+X�;
�#�Q��mq�-�<���D�7o}9�F2Z�L�NGp���v��XT07T4�Y>��P�n'�}�����%C--�����"�[���k��i�TUF�ޭ9g��>����!��ac�V�w�Re�4! ��n���7����Z@�pU��>�t���B��QZ:x	<_�ŗ�u�E�b�O�U~
88�S2.��a5���l�����#���%�31�M���Vx��J9�S��:�ȍ�����X@j8M�1~3���Q��;�j��s+�;���qpШ�*��ɮ�F�3g=^�Q~�]`.�~���H/�`��K?��}Ӱv�6������z7V&3��������y���dL��}Ϩ.�K�d���r�����.
ӞV1+���T3x�<I謓�ҎPz�,�V�枷�v�^��ڇ"���/{������V�����{�f̞~����ov��vI��u4ؙ1gU��U5��;�:cd��+Zx�۟Vd�\s9Z��ސܤ���g�X{������dR@O���^#ϯ�H��x]�?��mq9�3c ���'={J�9cVoo�c�q�n;m�����(�:�����y³�E2����#MҾ�Gsl�,0�V[��޻�	�Jo�W�����ag�K�D��~w����ˍx}�nվl�:��l��J*2�/f�p���'w�}T�E�TU(�����oҊ��$�]�x�������l��Hο�u�}0��F5v�K��^Q��)�	0�M�-���U{�܇��6�/Sqj���F-U�uY���ۮJ@���ߋϏo���2f�������k~G�����P�iB�'��J�և����y�M�����ڦr�����l�-MR7+�	��|�4��qT!�Ѣ��Fa����·&�J,�P.o'��i���a�Z%&���v�_�"-;/5|� jS}�j&��;��}S�u��*"��3t�.��|hY@�6#slpx�Lܖ��b�H:�k�} 8��q�ׂG:�&�.�0�Fɤ��E�5���c��:U�d�iF/v8mz(�b�"�� ��Z��4��wK?a&W��"�O��6]�n� y��(1��(�Bك�>�,���I䆥Yj����q�?Rrc�_K�r\�?�H�y���ʹv^b�c�UZ�ީ�]�;ua����B�xn��X��l��p*����؎���u{s� ����؆�����~�����}�޽�*�{,�+2<�[a7�,W�}.�|���E�/������`\t���,��87'��t�8 �CH�͟<�V�v(
�RQ�C�D~CE��H�Z/@7��xy�\�0�ʊ_`u�F���6�I9��A�pI�~�~D�\���dRRT�7?�T fڳ���� xA�F5�cG��,z� �_r+��{N
`�^��y[]��O�zP���^��F$J=D���y��g�hQ��G#2��H2�_K8Q��8K�$:���I�ڶ�Q⊘EoZ��~Ct��	�����E��v�o�5�L�\(t���@i����@���h�Y���ӿg�.��g�%������y��0�X���a����X;�7׊8ˑ-)
�#�@8�ƈ�J�����[ ����9����%�����:��
wvwA鵵��s��p�Ӆ���qừ8���<NH���gf��d��Ɗ&��ʮ88MV�����1�
�Xd�k���8���G�h,@�z]:l~@������ڿh���t����C)��P�qT�d���P���o�:(�%��fBSY�!��R]?o��)d�>Ƴ��S��0 �"@�E���WC�W���Vf�NN�muw�a���+ �L�.�nk�&�P_j��P���2j��d2�о�h���6.$���ՓEL޶\g[i�QFω�b���q�]Nz%F�崦�D�M�_�(�o31n���T �낵��@5�,6��KP��T:���8-�Y�z�Cf�U��=�u<���3��̬
m\��J�Iʖ�@�s]W�L�sA�Aw=)ޟ�u�:W�X��!]O=�N����C��K��X�j������1��3��kg�a���=�������i����n������-- ����]� �"�������,],�33w\13�I�ho���?� �{g��k��&��W�j���?�c�j�������3�ǂ3��F��l�g��ﾲ>5��(�PS��]�U;wc�5cU5�L2w\�h�f[J�����=���'r��&vI��k��&/��a���g4^~���%�k��L/�o��'��ׯ�A��f�i�$*a���=��s,��kgA����)��?
b��ӯ���'sz	�<	����z+H�mˡ?��X0�=
�Mt}���H�=�?��A�����%���j,��w7���77U㥢�B�m�FN}��=OE U���,��#�MxLd�=lE&�03���PXe��qt�1�(J��~Ԟ���!�>-?����e6���E!u���0��+��֟$����s�P&!5fG쬏\���c������ǈ�c�O�\i5���8P߸AWS�ydFe�-Ih���#���Z>�pwo���U�����2���w
�X���h����;�5�?�f~�Jg��;~yL����?8�^4$��ܶ��lk�ު��My��[��T��|H�}Q�8�x���=n^&�^�]D�ڎ�oӛVqqq���w�u�I�%_�ۢ�P|�rH�p�#��͏"G��v�xkg|�P'7&����F��`pqo2!0��_����J)4na�<��xǬzP��L �FvKm����a�
�f�%OAA`b�kq��_4��
���e�k���-���a^�ߥAz{
��DބP5��
\7$pbLLx��z�g?C�'⑼]-K��Q微ѯ�Tv5�����[yT�eǕe8�p�]����4�O�pIBb����R�S?l�7"՜���&�q�D�J>VJK�<+��,"m^^URR���K��ۍ�^�E��:99��!b�O���#l./���Dt��@��bFm*ی�O�=����zq�(-��,���Nb�(�`�\��y�? S�;�S��w댊UYіdSV�CE$ĕ�౯�Q_�~�O���ч��>>>�K�������\Q� 8ݭ�)K>/�	37Z��,>*���< Y2������Ԍ�w`M.���<$�Y-l�������EQֶI,ħ�BB���j��>LŹd��-o `*�q�c�-�j&�c�Lͬ7�iq�7�(���or����.?��/�V !�$��1���G��E}P�Xnvk?����y����h5��r�͹����gT7��G�R=��}>G��#���8d.F����i��y�� ���W���+�a����{���rN��b���t����I�J^ЇGB*�j�,�~$3�lm��.�VD}�z�}tf��9��_���mT7��L�snL�3,;nk�=��[M�g�����X����Р������M�l�^�Q��vW3���4��_9bs���ⓘ�G0���Ec��>�Xjs0ڼ���4��x3@ �,��2J,��3�uU���X�usʥ�-�������}rk����!�������'�6~�����X{~ 5��$t(���>\"y����R/.�U%.>��k����}���4/%p��K�k)e|�߀Q_M����������`��s�q}z��S�l<�+?>Pp:���у���>`��H����ZF�����=�ے�חZ��9����tN}�?]�W}\^:Y;HR�4o�����='��������Ϸ�����u^�B�p�K���s0;�m��O��]��,Uq���w�Js��2�5x�t�^�$
]� �``t�g���ʪz?T\T�۷01)	�Pc����~�$�B�Bg��
�[J�W�$���YM�����_}��5ջa?����(�1�m�_�Z�5���쇹��m��.����Cu	W�Ⲁ�wr�:�⪪�����t�_QP����?z�{������T�Km�U�x����t��n����k8�:�ܴ�^���C41�˥��cE��F�J��9py[�x�&��� �2���)]��	ڭ$;9�x2_��_��ߏ�vF}����}I\:w�q�za��"wW����_h���gfV�h��c����0��#w����#}�9L � �vf��â���u����O������E���т:ř�i�_+pt�5�i��� ���S(-`c��n)թ9ϻ[c��O�JK�\;KKeF���d���{��H��qdx��!�|�'��c�W�_zK��Q}�z:o�v"�}���de}�Y�~a� =��B�e?2�%+})a|�V8���U�}�.���h������	 � -�6~7�}⃚��v4�w�����h�L(��.H(4R�2�GSl�T�u&�VXH#�ۮ.2�)��j=oY�����;>��d�H���IJ��򄃠��ԥ��b���Pްq����5��4:�#��sU��%x��O�qP���v�1� �����)��'(��^X��O�	v[����	z��k���t���4s��u��a���1!���n�� q͡ݤx'@+�m}�(Z�LZE�����Q���N�5���Z�v/,�?��o:�z�����@��0�C8i���.fx��M������f��d���5���皠ݭ��[#|J�nf��
93b��^�V�^�Yе#�OD��E���z��`��f�Yqa�~�������n�ʍk+:��#z+��J��?�Aˡ�v�+H�`��9[��J@�Y����e�� 5�)�-ʜf/����S6k� �y�K�uӅ(�M`-��U�w)�X|W��7�����\
�����'���Ø>Ѷ�^3i�'�_<�º��5^g1V�?�]��9���v��W�s�� �������}�Dd��$N�� �z�h�F�w����%��*HN �������Y'�O�ͣ��z��R�8��2
g��(p��/gp�!#K=�u�}�q`YO��j��R�����+~�7qD$������b^���
�ǝw�����gtڑ?��E��������kgf��eM���d��������oN�mTAZ+�l�{�iq�O�ol���=(1&�$�v�G%J���!�n�h"_^cJ1��O)%����J�!����y��}�*�5)5��#��}T~�n�֖,��%S�4RH�_;e�˅V؊[���~���������*L��Ƕ�	�ܘ .�c��fzͯU5Ct��������a���H�5�]� ��u!���e̀���L�@��};9���L��%�϶U#�qE�~aCpf��7�W�~�O��C�8ʆ�k�[�`:��cލ���9����]��)9Y�-X� j�������㖛�/7��ܷ�y]�鎗�o�g�rGx_�f&RyT2�P+�s�Vlӳ�̟m�5��y�]���{�	���(_��ڔy��Ge�e����������4t�m�]�s*���)���䂅�Ӳ�+�z�F$���z/j@t�����Yo�E�	y8�xt��g���,�1ϻ4ZL�7:����q�7���<U���·�ʪ���y�z1��Ae Ѻu9��%��8n=s?fy-|Da5G_J�8�t�ك��pK�7�Q}3K���p|g[	�Zq��Z��}rw�q�����9�T"д�OA|'���§wπˎ�$�߻�(�9A���h�IZr�'����Y'J�yMe���lu��ғ��g�*��o 'F�?6�������l�=�����<Js`�Òk��f��ն��~!�z�|�n���:�3-��=s!�E=7�՚g��h�{�hz�+��s���anP@k��D�#$>��ɟ&��1�5K	9p�3v:��ܩ.��,J�0T�����(M\��#b3���b��W�d���.�X���W��ל�f7�~�	��"�����{�����8#*
���Q!��5��jv�YafP;���mu�5	b�6J�ޠ�*�wLA Ƽ���~C>����BJd{�}Y�=OL>5xL�қ������PS��˜C��i��0sn0b�H��y����]ɟ��ҳ�S��F#:���#�ݘ�/���n�R��[��w0����y�/���O�����A+����zn#/�ب��-��#��q@ }.5���+/��_���?8�5~�n��󊱼�y�߫56=>cd5(ii�1�b�7��~��?���W�8�Qo ��}8�H|�'���I=
�豲���($M�=����F�r���n�n*�kK-���6�oǼJP���a��[����[���!��'�/Do���5�R�K���G���4�,mU.%��"�#fW&�ؕ�������m��a�T^��<^U��ֹCZ�_4��K��YT�;t��m2�?By*i A(�[Z��۶Lʬm:il>t	��HX�}�?Tu~rq���yf�]ݶ��~���mN6���p���B���q�\<����5�����kj��Sj�M뺦�&�1�S����Ck�� O�I�����T
�~��0��4Xu%�O^�2�]V\b��z�,͆�i���	��7��ȊX=m��eM��
aaE���9M@��.��M`Yv��������y��{>�X^���~Uͼ��$�6FZ�9y�<ۈ
'Z�b(��OO\�f�MXiR��l_����]Z���{��-�I�����W��0�c�S��І�ʛ����� u�Y������BUz�=_�Y5Fx�f?�����?�Y������t6��nys�����F���sPL�v-���Z�@����JcZ�>'.����з�J��B�t���76ú���v&� ���
x��<E��t�@���z�_<˷+帴���]`܄ X|�x^�B��aQ���Ǭ�u�~�0��A>����4�=��׏�b�VV���y]\�Ng	J�[�'K��� �-���m1'�����y�)^���V��ˣ��ycP����f4Cִw����a���ο25�����}�Bv"��ݶU5$�	�G�������!�#�aK[�]����(�-�f�J���T�+\����EN�tu-Q`N���5�'�N7���}�.�}5�ƛal�B��h�쑁E �i���޴��f�y�ڶd>��.�,��vj]� ����W�����*���M?޻LusgQsf���[�K"�c���=�;x�;1��=�}t6\�=�\^[��/�����+�|<)��P?Zu�z��cO�#�ۙ�A������?U��s7� L��i��1M���tk}�8��I¶���X�9
���s���5��qHė|7.G��*H/������  �k�깒賈a�F�	i%�����c=2�?Z��'��qW�У)�� �x�1�{7�ׅڀ�D_�����NEq��x�8/G��/�,�3���k �cW�Ty��������ccFMi6���eŅU�N��eSݾ�>�EY	�J��T�K�w[-lo?�ޜ|�+�xzsw��X���^R��Te&�6��. �a�\��n�I�K���I�,veS�?y"B�١<u�������o��+��^B�W7�'�>�~��c��܏����S;�������n�!���:^�kS�hϪ�в��$���� >s�9�\��Dމ"
Lv��
�:��{H�ډ"��&�,�En��/�Ӌ���;���R�����ӥ�|*����ғn��>�(�h���yе�p�3{"خ�>(�}R�D��{��M�ns��9�uZ)��ۻ6�65���(�˧9>�D���RI��3�57����햃�B�s[~D-Z��Q<�^d��j�=I�X~&��V�4���t�κ�0�z�]�Cǥ��D矝�Wz���v�G8Ŏk�]Иa����q�o?B�mf�!�2�;��i'�>֏+��l'�(�q1'�>ѿ���ZH��!k_$B���ڃ���|�d�wzl,YUC���c4��,I�A��?�}Z=3���IY��H�r�r"�*ȴ�~��d�v	��h��ܜ��`�.c�������o�����mw��S-��EhM��+���\�$ca�t���>-���\��ee	���]v<�[k�`�G�� ђvC��D���a������]+G�L>���6q�#�����~����Q���=c8�׀��i�a5j���~/��󚫣Њ�,�,��*�և2����>�Y*�.��8I�>�lC��@��/�e,-h~��ZZR�a3zB�׷+�(cm���p�U��;���9���*��y�%x�Ĺ�>�B����Wu��
���^�� �PtTD��nG�d���x�LHH��\`*x�[�ɦ���?��꜋�?���儰�g*Q��<�M��|������n��W���s4)��U�0f��c����o?X�[����d����q|���'��8��������03�+�7��T���
&E^R*W�����9b"^)l�ؖ�b��?P K���z�C�Pz)	ksS�[��M�\2�P���'9�!�Gix�Һ�PK���Ѳ�2��/�e�j��5�^���D��g����'��j�P�6;��l�ZZ�Ex�H�w�^x�L�*HؙO^tP���x�P��Aitj�-�iV���c� f9ָbEV>�Fɍ�+��.�c~C�NL�D|��i偳��/0,�zڝ}�.x<�1D�q��0�UUU�穁���q�,q\���@(w[��{2 )���&9/�P*e�9G��b�
?ɡ�V�0�f��--p��S'���W�mٷ�ڑ�P�DK���`��P�C��~M����n�gn�y�"qvX}{��k���nnw� ��.�m�FU�q��-:#��	�f�g�4p��*%�^O� j�9�h��?ߩ���y{����+Y�`v݉eLB�&k�@���״�������#Au�<5�f�]��^L-;�]f�2�wRynW� !ִ��^�}	2BB K�*^��3��;��e�G��mwq�Uk��� 7'�Y�#���<�ݪ�rYY�õ�-3cM�� �������z�i�h���-}z�ɽ�+rҕ��XTܮ��}��u��x�~�`��5w!X��U��~n�j�ZH�$o����Lr	kZ�*/�y/��A����A��C����'7�
�E��r���c,Rp&�Ut����@�v����>��ǲr��c;��'��(�7�U���Ը5: _Jt�K�����F����թ�5ZB�[��k��\ǭT��Y��쾙�}W�AX�!�"�'8�O����Xmv=�������b�����q5��D���@�0鏾t*�,�ua�����Zp�[�K�,G���� hq�&B�oUe�쇏b���89�W�\��A�o���m<u<<�=�.S�(�ۈ(	q�$���'��(t�z��pN�3���\��:[�I�j�R�4���0�7���k_4�U١CYiuD�Ղ��z
>�1l����?��-V��=F�Z�H�����z����L-	k���S~v�Gcn;T���7�s�q�I��Y����j��WT ����q�]B���1177��Y>���D~����g���6����d	['
`��3�����1�l7�'�*z���4�"�)��=�]Ȯ��3����bt� �O���s8�wQ�&���B0#�[E�l�`��Ǻ���m�S�	y�h�wHJ�I�I�l����Or�NQ�(��[R���"r� s�N�T}���ir!�a��Аl��s���!m�/�u��g�g]Wu=�!�; �r�Fz��͇�R���ւ{z4�z���4 ��VE�Uh��*-��� 0�C�O�I���2ǣ��������JN�w�QX%ʻo2E�>CHR�&�wn��l�IڀKCI���!,u�o�r��#�Ԩ6ɩ����ǯ{ο�7��#	���v^ty 钕��0}�%D�ݹx%uyo�zG��'�����?�����6<X`-�G]r=�H��f�/$#"B�m.�A�<iii)�
�x�>޲�����X
B�dB��S�>f�8�Q_P�T}�B��{�r����[��o�6B��2��b��rr������R�NGRS���S|��];Vn� &�'$]�8:�;�fw��9�M��3�/}��Z�z��i�����'D����(�C+6z�9���@�(s���Xb��?�'����zmc�*�P�I>g��/��99��/(
h����0I��7�Y�;F쭓~�ϗB-(*p�s�T2�L�Iۡ��&��n�D*b�>�>���a�*>���D
E�U����~8��"����[����(�":{���1���{L��*m��X%�px�q���i��o��"
�cza�~�(���	  B�*��-��^�=��^q�o��7
�G}������ܽ��4��L��4���%�,��Y0��i����R�d�g���-	a�]�S�j�K��7�(���J�"��ɟ�>���z��w�
~�y��..^��,��DA���e���AB��a�x.D��A��vP�C���c=�$y��[7�e���	�롴������v�dd"�9"6���2���5���r��I���6 ��>�U�j�$L��=_�w��1_�L��x��YȣW�΋���q�#������}՚+��W����
,����{�y^�.	^�����>�/4DZI�r���e��gj��������Θd�	�t� ]�Kb�хI�Z.I��1��0ځ$�} ���Ā^׵C��a��� �{}�ߵ����l�ٯ̓4�+!*9Z�Ɂ�Q�NK�����ү��F
�#h#("�S�O�ko��YK}��b��y�t�\ۉ:=��Ca��K��0�2�*��|���\~JH���ʚ�&H->~K�'-Y�=(���OQA��!
�`�/� d�Yי�̭�"o���J\�_� �!���{7��o5;��zd"z�P�^��v�-XL�(l�Fcj��1���!!KTҤ\�d>���3�SP7��P���	}>�P���& �ߛ��B�t���Xo����n��ɇ���i�9�7���R���y'K��k�����9�	��j�����2��4���2ώ�p�ܲ��5����ʹRpB\^����l��f�F��N��*���>�
$���qY�W,������2Y5d�e/��+�f��n�� �13v�O.�l(��Y���'�����`;!��v�~���S��g�f���|*�8A�c������_�2JDc�͆�������"X��!�o��vb���ѝP�WP�n!�L��?��qCʔ��$y��ǵ�ۑ���/@��ګA^	27$/���m��(߇�t<�h���We[���s-����q���***��,+"b�s����5��u�Sܔ�����j�;{\�ex�~P��9y$Aә�=8=��	����,D�),��qzگ�
���������ʿܦO�ka0�6�ǉ�ʼ�<N;=�O�}vQgE
g�͏��
�k����:ߩ$tTw���Ѓ]�B�^�ƃ����ח�?������jc��9�8��f�I����u� B��d���*���٣�s⻺��[:^��*=�˼y�!p����zF�vޛ� 	����C�}O}`��C���a|ś��婯���p7�C����J��I��ہ���Z����܉tK,~>+�c-�Z���#F3��Nq?��<,JU���Ԫ�lw�w*�=G\
%����7�5�iS6vv����Q�0h���'h�����
��z�j��Y m`9q9������b�(�$ `S;��Ӏ�$-��>4���ݝ���@$�[�-��C�\����VC���-��Χ<�����7�|�E"��Hز���99:��u��B�2gO�D���us���#���
T��.��U�X!����
O
�e���
��RC������������r�o"�g>��ԛQ�~���F��X�6s����/�{Z�33��0E���g�.*��#�&���$@a}��,�����+9��Z�T���jʞ�H_�<t�~���RY�I,~��e��M��D{}�҆EBK�����S�N��T�l�+�X�	��������		���q^͞�/گ��bB�D%)D�M �a����x������A���4�7MA@�ī�G������fu��iۖ	��]""44hw��A�E��j��,dhHT6>��O��T�z3jdo:w�{�Q�/��L!����b�}�r���������h�@D��C2��N�����@�X�I.S��Đ�%*��sD����X&]h��ȳ$&��l�~�p��ԧ�c��2���)1��6lD�}馋��J�6o���I�V��`���٧�]U`�W1�J-֠h\���̓8�\�,i���R�E�����ô^EOu��3�	7-6z��In�4M�"�
�.�4]R :�����Dv�������eM�q�0�A д�sɊ�Ռ��" ���?d"�PWȚ.%�����=��OG��T��^�B�y���Wf����ن�D�<uBB)��!��&_S�W��h���Y2�w����C-�訠UN�Eӹ1���%�,ߔ��ڭ���V(,�/{,p�ZA6�;D6�V�X�v,��  7��|L��<0�tBV�w�ɲ̐w�-�aT��vw�F��q����G���63�Te��"~`B���Ԙ;?3�_��[�`��>f��!��.j����&&D[D����l�NY�Z��\\�xa���n#RA�U��É+x~��\M
��&�<�T������g8睿�s	/ M�+4@��|o`P~��}⯙�����F�:F㹊����O�cWA#�?�<.�'���\�թ����UH�0ek�[E����\%y��-����I��m'�gm�b�F���D��e;���*+=<�?EHr������������\���Vf�x����m�i���=��˘���3�[��pp�[+%���D'���v�+�ǝ#�+UB2���M�0 �̝��b��P!A�0KH��Jc��o��Cr*�2�%d���g�[�F&f{��+����~#��L0�|Keg�^�Y���d���T��Bk+����ԧ��Xk�"�^BA���C�k՛u)c$�Q%��!���7�cE��*ʾ���o ���
ԁ�ځ��Y���L�Q��5_y���H�#�̻�u%�J����@�*/�R�R�����nntw�����b��I./&,��ǆ]>zdd�_%:$םa쐮-R��Mj�� ��2�/������Z�I?K���r�zh��?�|�RҊU,wI�Ӌ�?%.��è�(�!�,,v��f��	
n`ȉ����X��l��t��	��ּ�\K�A��_hםe4�e"����ޥoj
%��U�avV���1�P_b ���Id�:sBa�s*���+ܦ��.���L�;��<�Xr;"�/Ύ��~��c���7\q���B��z�Lu{��u�#�Ȼ#��d\�*.�u���䯒��4Kj��2	@TDY�ʬ����)�l�ԽC�:yڡG�����X��1l���~
�%u�Yg�+	�s@[W��ә���fMٮK���
�o����?&"�k;�n��9�B[Y k�N�k���������e�6���Jq�/�\.JnD�"��yt���1�e� Hw%}�;,d��@,���4�3����r����?*z�z �{-�B��FBC�9nh�� t�?!�����*�{�
_�N��/e���>�n�`�ͺ8�4,�8�4A�b��÷�I�A�'O��qg��櫪nx���ų�P���	���Qm��隴�b���,C����{�>�� [�L5t���-Z���&�Sd)g<Ā ʐ��PDQ@κjUe�<:��dFl.���by�%(���nGKKU�zqbGdg��bWۍ��i�#ԂQl�����i��$dee������JGF�a����c�-Iu��V<_1y�&��HC�O/�^H��s�3�V��8'9��&��CM�O!��_6;5 �'��X3J��+���{6!,>?��l��9Oprr�J*���(0�>��jB�<��ʉ�d���bL�v�`T�_Fbak��)���{�/$@�s�WJ1U���٧����W���
(���ؗ�ׇ��ř0�9�x
Ԙ�jc��-���I似xr���k�������k_0sh�h(�4i�ǮR~�
��~�(Y��� �f
�d���Y���*��d������deF߁*�� �z��� �a��c����u�	^��O��|��.�x�L x�9�ז�*�9A�9!s��%����܈gZ���@7�%��r'���T��[������zWJ�K/<��ˉ�~k��Q6�������j%�vd4��e^�-�i�g��@��A����7�л%4���P��ͯ�������&Y���G��)����(]�����n�K2?h$�����O������G��\�&&��U�y F[O�U������f����b�����l���͖��̞�zQ�	H ���LI�Ҁe�N�JHԵ�F������h}���|l4_E4I\PP@=��zvs�<��N�_���+.�zC?
���W�|yt͌GGW�J��C���>�\������-��~�ej!�w#�#+Y&/��B'�M����E�^�/!�M%3�\��#aH	�	�����-��-�k�wW_ +����1z�;�r���!�w�����j4Mbb���?J��]��P
W�&�$�� ��Y0�z�Y��܃=IkQ�X�NO����6���ʂ�!��?Xg�X�����Hgrb���h�=�d<�e����{ɧ�Ut?�dͪ�@A��Z��K�����/�99�2H��/+c�T� 2���x����26t�="ڧz�����~K�R�[ZaȘA*P��b���2��{L��N�Q�L�lPA����3�u�Uw`l0�wi��"P+f����P�_^\�ʗB������Ip_4�8�����G�y �xC����!�$UE[�}sK2�/��3�*<DdRoUk��D������ �����#W~�h@�9[�����0R8|B�5�p����&D��lS4��c_��|}]��B��3�J����N8f�ma2��r����8�Ϫ�����F�]�#��2�XQ�~���`Ԅm��E���!����7w�W��{�k�͸��!�������*]f�{}� z6p��:�|PQǂ�����Ժe���MK��h�3�qC�%q�����J��lYJ5��d$~�H ��}"`� ������L��\=�؉�-�8(�g%o�c�P�㭖�"��+]��C�N4(�oT��iVP_d<�>J>���[�As�r��!h���'X/�J1��_9L�W>8��8?���˯��^ޜ��N�B��v�7���V�^� G�L�)�ǆ��q�!��K�	��IA#os�{���<.�t����:))z�f\_nkP���"�(|����Η ����iX�Kǜ�Q�� d����Ū�Pƽ���9�)&��m�s}�V.��^���
x����@���[�&s����/Ɣ�W����]��U���5��ʝ!z���V@k�څ��c0cښ�G��뼿���G"���Z'?��Q���oή�Vz2�� ��\��U�t^�r|87o9}���VQ@5+4p�Hp���a/v�Y�Ɉ.� ����nY�؜��ƓV��������6�,M�H+)�9v������Sʴm�O�@Q"��+5�2�C*���������@8���C,Z�/.�)�²nO�Iﶵ�S����r7ͧx�(U��he��?\s�v�*'�T'feEѩ�赻*T�`a崴�W����?K��58��@΄��K��Ӕ*�<���FW�2$�&����V�)	�.����3iC�K�-���q?hN������|�HV�:��+<X88܋�Y��~uuu����-�+M�����=Z`Ei�@�_��2����c�,�K�X�J4��*��� �5�y6�P���nH�t>!��\�(K��ϗ����+F6���MJG��pu?����9�T����Qi8-�)���
h���̴n�w	ߤ	N�D 5 Da���5dhIc̲]�L���ߺ���J�
�� ��݌7��S_ƭ��
޺�B }�Ωծw�v*�E�uCAN>��q�X���`�6���R��_����ߠ��O�BN� ����ƆN�[��g�ˍb��@���Ы�2�t+�p/���=��%����B����=nB�=<���̨���5�����"-(��^nb���]rM�`��Iȗa.� �����E�����1�g	5��s�Ug:GH.�zB&�a�7�Br����)��2���{C=�11�{JE��m�E�=�F��F`�~2�f�g�T�tT�b�~������������U�A��s������ֈfuQ������C���7���֠�o�o)�0�G��$�D���U�3� ���U�y�׺��q?�ZVK�@wZ�L���B1i� i�P����SQ�ĕ��L>Z�����V^��cC�~|m��$>�>����2>9$`�%�s=N��~{-!�����W"���[c��+�^�Q�/Y��׀�ݛ�w8(-�5a��WRT�tw�EU��n���p�����#��@�!4�\�����!n$~s��ۀGY���- ��L�؆�����te���/B��la{��>�oų�i��E�EQ����SA��'H�5�(��I �F �y�v=2�\}K�#�E��]���:�J����3oxnJ�n�=�e����I�E����]�r����������g5_����@)3E�x���وd�=?}�<�E��[�IM�{����{L��-����eh �lv��q�ϡ��%�[���֫F= ���e�d�Ӷ�����ʿ����TEC����.M'��:3$D�f5F���'�j!%з��mM�9ˊo�e3��'���A_Ƅ�����Vɳ�귔�����q�Ci��*��x~�AHsI[[f��#v�0(i�lA��>��%���b'�H��Â�%
B�R1���]�?K���)�dǗt�ޠGV �&��)|�!mA6C���!���TF���&�Ř���*���!wY����]BF��o�[)�#q����?ι��Һu�QN?�L�!������v�CuwY6�TN�g<��n]P�H�������E�R
�<IY� :��=\є�V>���T38�&��gG>k1%� iR�@�a�d(��^�&5@@��*��B	�e�.�t���V�8yv��U1���pY�H^���v��c�$���O׈��h��������d�2l��	�+x�U�ק>��V�8��f߆1��Y�8GPY�NB���E�I��:6�#��R���W�NMM�w�0IHLD^rr0�D�]���Ɂ��L]s�i������͉^3��g|Y��"�&21R��ڬ/�D~�VU�#�b�����ck�ħE�Z����N��c6�.�z:g* H�<���?��s����U���22��	��w�8��CR���<Ѻ�;8���F�(E^:뽾<1�$�8�߉��C�m�L�D�2�bQ�˝��w��R�h�������h�ڈ$Pa��"QMHJ2����0cK�Uo����-2eO�
v�Q��
h(�rϭ���`NƷ�}AU�Γ�n �IH���w��X"�)�a��c�G�C<�v�����d�t:�|P�\N���c
�����▇�����a��˨(P�u��3e mg>���Z���5�\�.��d��U��E�А���0P�DH��̪v]*�䲔���晥�!y߻U71%*�?�_�#��������#Rd��� �dccs���dԓչw:�Kx�x_У�Y�M���t�����0���	���y+�m\����,�P
˕´�?�U����x���٧y�SX�7�{M;24���1�9�X�k��UU{��׭�आ�0-�w ����d����_��G�`тON�9��$�6^�s&�.w��pT���'dDl�s̟Wj��"rY�W�[����ښ�f���r8�7� �}n^�b#^,h-uMC�g!����������Hn�y>_�
�Giq,���ua�)�|��S�ǥ�J�>7J��9Y�2�uKx��F�����n�����5��X
+.'H=����E�ֶ��,�3� ��~%��[KP�b�/�؅�77��"�q������>,'��X��4��s���H ��	�����U���6%�� ��b�=��nd�a��V���1I���[ɀ�u�L3#Xz��a����Q�,�**$@����A{�zi99FIg��
��-�-?x�b�2<7ư���frk]���Ѓoʓ> ���L���5�4sNOO�ZNQ^Σ�=up��W�	`���]Ɍ'���)<�@a��lCOdC������!.惏����B� o٠k��'��)�@Fq���Yzq�#���(�o~s:�	���L�7t
��@��y#�P`�|�j��]�C�����/����_|����A�X��M=�V��B&��rY� �~��B�ۿG̰�!�tǨ��6���ʤY�g�+
���D�ju�1â�1(����?]�_SSs����BDYYٴ1O�.������z��= ��ȷ��Rb���V�ƤH�Jk�����w:��y��fryHe���������H[<��iM�@�8�2�h19%�M�'G��|��(|}�o����N�GW���p�9�I�J������0�5)#>���x}�i�YI��ڎbfd��y�5��T������9�����С<Y�
� c
Q�/��ܝ<��G�%!�f999m��ulll�O�,uz����n$��hnl��/1���+�p0)�9�ׇ���GT_>����&w5U~������yD����]�<n�f�_{_����?T�B"B(�R��c+["K�([BvY����^�,S	1��c�(C���G����������^�>��5�3Ϲ�}���z��<���[ڛbNy)H�q7���vhg��L��NN�߬t����p�.��_�wD�:��j-n^Q������7�l�]�d��TVI��UX�="(r��D`cY\� ��
��G�W�DA����c��ݿ�� D����(�� _C������`��+���o�zѯ#]ëL>y�-��. ��"&��w[0���
�o�g𴇂��38��7�'�o�{���M5��=��j�YP�'���I�� 5|k����	q8~���U�##����楎��v����1|�_�&	
�˱˻5P�]T{���c*`�gW�ܾx�q���ل�D�P��CƐ �iLzD?�jsz凅���]Y�!�Z��g`a1��)��S�;w�Ɛ"p�Ѻ�X����3PG3�R)�9?BN뗘%�l��Do2���7/�q�������5�m���Y�ܽy���(Y�?7��U���V�#��NM֜�B+^���MC�����u���,W	j�l�]�n~!T;������Rt�D�˗^lɂdѾ��!X3�.�늘�b(\>��1xd��%bP�}���cEw��@�����X������Y ��ŝ�ΐ�`�Q�S54@?��oe�����h��m�B[-sO�rso�G!��n������[[^�'��G,����>�Dj�������0���
Eq�f��H�������L��A�|����>���=	"�|���������[��
��;�܊��r��=��˃��3@�b>w<y6���uɁ	����Ȼ��dl�B�Ĥ�����"�ٕnʩ���-9��l�G��h�����f����A�-�E�:����.f��L�S|�!k5�b��V�~Ŝ�u^R��^pd�@+8���l\(�v�º��Z�P:WO1A;ņRO%��_��J�q���:qF�����ݭ�WcÀ-��]d�e�~eB��KyR,���3��<}Vˇ��@R �}}*I�oZ�(��``��� xA�%���f�J׽+g�����h4����M�:x����ҋ��\��G��i߶��^d�>!i�������~��rY0�[�ͼ�#~�b�P��C5�����(���oQ~|#�qGe]5_�_��3ϸS��oO�t�~ݙ=^p8�1�eXpS(q[v*���~�ңRO��bF��@(��q�)�)��Jw�\ۮ){O:$ ���ҏ�Ykj}���j�������pj�oTaH��[:0�6OW�%;��]���0d����^��y��b�����"ۭB9�4���uqHe h&�s��I�2]�4h�U>�&�}��}#�QU�$Uj�{���n��iv��HSh��#�!<d>
�,Ӗ�=��������tˡT@V3]�pa��7�����Hd{;�+�}u�DXF�|�_����ǒ-���GN\��r;�Hb+5,^J����D���D9&*�������1�Q�'41$��Ͱ�ZLs/Q���;w�&Q��������_�U\72J���#���=]�M����WX!j�p�T��v!c\�������%��Z�wn���5G?�mi��}��$t�m�.�GDH������4w��w��6�����5�7���c~Z���:�$s�@���d8� M{fyX;��晡����JI�t���@FX��m͝��?%Ư9���#tdZS�|� �����Ҹ||���ś��$���騵g�1C�	tn��� ⍘��NP�T�xQK<�
��F7��0}|����c�'9�D20*Y��v͕+��-��i�o�Y�
��U�ɑRZ@��5
"h�稪�Ў����8.N����V.��7�;��c�1Yr��N��:���L	���p��9�uBV���E�̋��#�n��NCB�����ˡI��Zq�"�.5���2r˨���
�B���t��2V�k���=���23���߿I��?>Y��E����ԲxVˆ[��/?a/
5�Nt{vgO���@^#�̓���������mufĻ�E���<I&�Ύ�����7�t��H`FOO�b5�����vV�vV��� 2O��8I|�0�.�ՠX7ޛ��3�r�0�����cCA� 	#��ft��K����I9�����{Ɵ�6�d��E2}��U&�����/�͵j�?_L�O�����} l��j�6����ۧ���?��@�88��RK��0�����F�1OO��&{��o�]l �!�
�`N�b�ӎb5G��\<'>���g��UkHT�zA��1�����&�|��Eٌ;�pC�����/\�����R�/�v�-���,�R�,oo1K�R`�#P���]Q�w&0��
,<j<�7�* ���>u���-�&�����9��4"��-���6?b[mS�#���ۖ999���АEW(	_��<s�(��������Z^�u��ɧ=�}��d�ә;SI�{3:��Ѱ[F�z�~I{���_=�x�s��h����g��;�[��Re����H�5#�dч����M�	�o�,AmUt�A|JJ^�T��R�HC �8�.��q0l(z/(M�rO�\y��5&��X&ۿ�E��r�?�|ǐ
�4��ȕ���k�$v���P��ܠ�D(�C.��Ί�xg_n�d�~���C�3��z'm�������b����5���NQ�H =�C��s��f��:���0v�앾��N=��!����1(�XJS[���2Yq����׌�Y��!;2����v��4� R���ul��~�F�,Z����!�'z�%���"��@�E6
S@��?�~:���qΐ�����ŌR�h�����Z=�,����4o����}��#�H��~��Y��c��h��J7��K��b2BE�V����a�z��7���	^�ř�G�XG���	�Ꙡ��ϟ����˕)��|�"l�FOZhv)$�@Ba�s/~G�{h><-�����R��/���y��4p�2p���W�p+	�ґ7z�
��!�$3�m�A���x��_���� �Y�/���x7����S.M8]���>�=cip�*[ �i�p�i9Z�FW�5��/��V��=N�e���GBu���g�9)�k���,�u�O��;9??����"���Z²���=���<y�[�p�C����aw}XB��'�vY�)n�\���V�=1���t7]FS.$}r[���ԡ��w1�����2%��￉�e�����#_��b��z�qP�QNUé�1�54�
�~���ˇ������]M����h�Y�U������b_3����˘��A��'$#j?��	���6�u��ih)
�2tKXq�;��#z�.���?�UK���D�Ӄ��O(@�蔈�M��W'B(G �ؑ�3�g��>����`����o��a�POD��-`)iiPݾn��#��nTR���,�6+>9�bqc�L*~˶�u^T�8�ų���������a�gA�iM�O�;q�'�ď@+v�0H�|�Pd��+�>C�ĭ��H|\��[�q���
?p�+|�ՅR��<�iD�&����&���h-u���x��֛ЍI�<�����!���{�D�P���h�R���4�
��&CS��3�B
\2�$:#�����T�ϩ�M��KK��۩v�u6�)� ib��Te.�P��G2�_�[Q{��S���x<$��?�����x.�`T{�t�r����ײ��"��]�x�{��V�*��H�Ę�/��6/]�ї ��47~K���^Y���1��ɽwZ$��Y����Xm%���c�nZ��B���g2kؙ��ʐ��7L��eHJ��d{
*�{�?�e�3j".< 6��>s�N"��f�o��
L����7��uf����%��?��)��������A�����j-�q�a�K�<���AwP�-'�G�0Y?��ohbB�ahUn��������n������P��EЩɡ��P��>�I��U��d7�y)�d�L�����c5�j���ʖ6���**�`�c���ڇ��qA�n��Y^|�W��b�F3xr��.p'�ؕ~|P�*"*�&qF����Im��&�P���'��S���x����ٗ���[����#�0�oߪ�ݖ�j}t=E�*p�R����b��@5�LtlO-Q�K�λ�����\����&�����$�?�1v7c������Ɵ1�^�'�)��%�>�$[�t����>`(V޼<e)�����T��7l�Lv��VlV�m��'�D���F|rr��D��aF� =��y�:��ʈ�WF�$r2�r>����?�^�����?���|���No�e���G�>@Yc���ĎNN,LQ֕c	))Q++� QCN7������U�+�ru�X�,��*��V�W.�z��E�1���\�#�XŒ���Y��.^P��N/�8�p�3�N;)GGǓP�df���)�B̆!=��X�:���yu��_<�w�ށ�������-�5����9��O�?w�]n��r�|���|'�BcQc����@bB����1�0���J&=!--�LL��=S�׸��v�I�5����Q8���%ݏ>�KtV�gq?� �����h'���{L�w��֙����2F�s�Z���`o�ύ���306�C��Իv�Z�c��JJ<�4�q8�!x��5aC�$V&�L�>����vS�oڌ�����j�f4oC�۷/���o�)�E6��{t �X�_�,#�ǡp���poɺ�,�ŒI����a�0�<V�ϟS
��;מ�����&���`4����)���T�S0���Y���s����]�m9Y�3��c!��ov8z���PP��R��.C�[�n1�o-��^>�Z���h�
 B�޽a����`ur�����t.���OE_�gT`�6L�Zl�7���
6�ď�x��2��_�%��N��n�Y�������"�z
���x-P��F]~�@<D}����C!���4�#Z0&��K^�R�\~�� ���4|,V�<�P��q��_��ץ��QvR���㫝�@�mlx�91�Vr322� �`'�ڃ&�<�����]�`�[�;�������2 �_2;x�ԏ�*.�2���=!�^W<��(�e������q�h֜'�m��Z�#�Zg=�K��(������Q����M���.�Կ��H���[O�b4+**z���[���'0�h��;�x��`��n����L�� ���mr@^_����=#���K�?�q�P�|."�-���Z!�~��������<(��ߔB��hol���H8�~^�9��.�Ծ{�7G���^�jc�1��p��reM2�����'s��y/,�������`
ބO>P.B1�b�ӄ5�ia��\|�Or�ۅ�T�?�H��0F�(��yue)������x�IJ2����T��U��8��p�?�K<�sqk�|�K��޾�:�{��p�8nq�׬l�T�'F>zPj_�G'b)zHxq"�?x4!@���H�c�&o���Z㑑�џ?�Qy�2R��)�Zqv��b�MS����ʎڼ�+s:)���9��#?��Y�p��%�<�w�����W�Gh��R��6�����`�}G}a��G�eoW	���=�wѴx}�W�9���4�j���Z�I����>���Ƣ�_���s,7SȌU3Sr�6�+I���-�|��3/%}��^��Xhs���6+4~��KNNv�ep��1���3M�J��dA�#T�qh��`�����s��|�����V�p`yXp�"�jTJ�f�k�y|�H@=;�;N����񠞴��i��]�k��z�is�N8��ᢥ�Y���i\-���M�x�1�����1B�7���M�G�ʖ{�yn����b�W�M�sR�T�O�����������d���.��q�x����nF�r��ڴb�^�wC�f[t�r̈́��E]�'����f�N�s�g�[iҏ����{�vnM�<��<�ő�����!��ݳ[�2���2r���&����7��/(>�Hc�ͻ��[�Y�fYU|�V�ȵ_gC6�U��+����X�n�^������Wg��(�s{-�k���7�1���?~"x��e嫮�{s�>�T>s_��<y�Veؓ6�����<���$����*/��_�jl8_u�v�4͜w���]�QA�O�R�����9�.��'R����0�t�M�8�-:#�s������:Q�|wO��������.9�4h���H(ľ�q�YN�?^����t��#�C���"nnãa7
���P��z?��Л]e�����=�|�4�2y\|n��Ӏ�_0�N j����}b2C���>�
���� '�x������͎�Ŋ��^��jK��x����:c.{���OQ�\g�0^���;�m����� �8���+m���V.�5�4�C��T�Ⴌ�G��aT��~dw���Ĉ�$�W/*>�&�ߔ߬�����{as2�y� ��ss��./?;2�2[��7HWy}��VLQQ�B+�e�|�=��3�<�̟�����9ԡ��uh���*m!�@�Bԁ����r~n�$�g{_�2�!U�����d�����d�	�ZX�w<a:�|~ߟ7L&FG/�؂9lÝ��l# �6]�����:j�G�J��d��yQK����N��Ok�Z��zgw���LN�3E�vp�G�l� em�Wxz>*�Bvw�?�/��}�rx.����R��.ܓ
y:�nJ�^����ё9T��b��-�=���Xt99�E�Ȅ(o%�m����U��u�6q�{�(lD���L]�O�o�+iŞ�����s,������:�ܪ��`����Dc૝�fW0��QK��{}Ŭ��';6�ڑ�	l}��Zc�G��|*�&�Y�?��p.��x��A6�t����Gi�Gd=u�V�p�S�[̖����A�:99�����]M�|��?-3o���#vv�;wi��[S6v�z�2�Z��tm(�������92v��I<������(�iF: O}G,߯a���u��3�9:)%���V����٤�$?����L���l����:Q3�֦)fِ�ݯ(�M��(g�����i�鿶��7˃U�,/��:N���{AI]��Xg6AKr��e�+B�+�c����}B�R��f�l%�|6.���$���\�r���[�eڽS��$�,1��bc�N�obe����*�L�r�..�Y%^*O/g�����������m@ �p���C��.z�?��?��p��A&C����:����l�I��&��Qz&��?�"�R!�&���ŶwQBl,F��פT�T�Ȭ�E�� =@��K���ډ����y�P¶��C�5���mŒ��Z2p�/}^!���-fWP�~Z�O�9uJK5�\LR�eo[�� e������Z	���`�"��d�\�|��f��1��ܙ�?|8���hl7�/!!�������VAe��EΪ�k阳
^"���<������(��1�O ��.��J���tX7H�`/QR�\��C�����G��o���H�k޷��d<�u~o��U���b�[H[Q�����
0uq�	���KK�K��vvv�	_{''�q�. 4�SR�l�B�Q�����i�ζ777K{6��|pM%mow�P¨:����g}�\٫	��J1Ⅾ�WY�>X�=w/7�}�F���ؘ��9���[@;�k���t����EEE��jօƢǏ7��&~�M��9���4��	�	�B��!g�ݵ鲱պ�Q'�3� i"L~˧��d?00Ѓ�����w�ƕ�@�i�hf_\[q�����֧�UV}������K� {��hqP�N��,FW}�H."�;�з*�N���2[�0E����@�n���t���>� ��E�\��9�?>�p��RR�R|�&2�J!���p��|h9����pm��r�B3���6(H)��J� �;{�1ff��f��U)Ga�F Qa;�4���f�2	��`. �iB��uE#�E({))�l�K���Xu,��N\��)�9�C�����TT$[�d�޵�Y
N N������Ya��@�g��k-��C@p�^ ���ǧ��!��8���NFq�|���/"�k���)�i:֌��j�����z�G�����i%�쐑��t�=i��-$,<�	�j�حŗ�l��� .���/z�;!W��E"���{�vę�s,Py���A�����1k���B��,�!22:��[XXФ-Ү�i%��%����peee|%�3\:���[�YZV� �&?A��>�߮u�;�}rM߯0<?���6�jpvs�6�<>Tb��x��ݻ�fCu!�&�0X�X;�C�����V��&���l%q�r�6���58h�P-�ǫ�@t���8�����:�#�,���APC���![��W�+�
M�ژ�Z���|���/ �V/���h���yߐ�M/p��ʤ�$�����]ͯ�Lc(\��Q׷�rnmx��`�9��z��5�8T0�̉I��&+w��{fFF � �4	ͭ���Q:������
U����j�w2B*�|�4{6��| ���%G]�p\!��:��@	w��h6 29�/Gz�vQ���K���i�zx��SD��}�I(����Qu��_�����������q̊��[G|�{�a�ecW��9t0^��n�����Zc���$ѴLcL�`�� ;�����6V���bLOh<�y������{`�A��������ެ�*}��t�u%\
�5�j����!�cxkKş�}���V;� ��j��-�A���W۹�#��7P���RcE}w�A�5�ԋnX=�?PK   Q�?X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   �?XLe�� b� /   images/d88fff2f-2870-420d-8277-ad43f3d18502.png�eT�Ͷ.ڍ6��޸�5.AA�C#���@� �!H�	�]4�]� �N�Z{��=��_w��c���oU�zf�YSፅ��aSc  <ue}  H
 ��0�3opu��_��O������=��\`���0F���= � �.�2��:�%Z��SG��I�Bg���{J����]^��ѣ�pR�L�Ě(��VgWʝLs���Y�ʝ`'%�	K۔���	�L�s-�1�Q9��o�K�$
?�L��zv2Z�PN�ӝ�2O�&2�_ٚ�_���6c��,��7`����+����]d�o�i�:%��2_���r�2 e�rRR�j()��HHAr^&˪�BI#uJ��Хc@|**�O��
�L}��L3ixx����?�<�3���q'C�f t��P��<�(�`�ys�"}u��)TtT���F���b�W��@"Q�@���P����?�#��Md5W����B�51��b���r1oY#�s�{
p��=�}o�&�C�^k�H�P�!_4v�}&�t�i���E���3	7�g��3m!�ռe�u�A<̡��ClPa�1U�6�*;����)O�g1(%�b��?v�gE~��D��t��%�$d�C}7�N�Q�LG-?���Ϛ�^�v�1���g�a�Pu[�����H��n�^��v��-���s|�D���I�Y��?����ռ�w� �Y�K-�3VH��uB�������������w�����w��u�y3���\e���t23:��2�jh�+���=a�:Om�m%���e��� p��5�?���K�_��o\)��_��̌�x;�2kC��<a�"|"|�*�N�B�r،2�v�R�ʪ��@�d���ݥ����������<�%%%�����x��^������^,A�C�e���������������[�����_烻kk�7���?������;� � ?���;��U|���;��"}�_����iS�z��+����w��t�[;[~��$�Bb�K5m迩��	���.�����������V�>��C���$��#)e7[�����,��);7[';����ll�DĄx�`�v�"���ֶ"��6��"Bb"�6�������m�j�
9��āYK
�$Dya6�0^;�-����=���L���f'.�/��NH��v��S�e�������������H�`��6b��b�6�ւ6��v��C��J��y­����v��:���¥���B|�3u���Gn@���������,=u�����ҧ�����������������=�yz!m�/TA>���u1������U���SJ�f�������E��/ƿv���6ҡ쬽����aHP!)A)a����R""R�b�ȡ��л�9��Q��>�2�P������S��)��?F��8�c���[HY��C/k_��-�:Z�:�������w��ׅKZ��
		��HJ��J�������K
��	�
�[�;�������'L��G���V������*���s���C	�����qf�
�����������	1E.��.d$���P�O}������0���0���0�����`�O3sEV@~�V驸�,��°y���w��Q����rW7� �{���}�CNbzkh�`�y$��� � e�����0�@�����f���>F~�od�9"�q1�@�G{Ә�JN�!�����C�v���EVPu]Q� UА��-0.,0�֝������^�AՋ~7��V�g:r�~�.�9�,)���:��4s+w|.�/P��l�I=�2 ���>��+��?����/36$��78��1BH �;bԺ�D�297,pb�I&�N9�!���GL����Iy�A��`�;�!kѯ
�!׽$طǿ������]�嗟���O?Wk>:ѽ�H�ҹ�/N#)��TSR��A<�12�4BO���x:��DOqDqL��߻y�n_q�^�1d�<�������}���L�W�>>8t_�송�]������Η���:ykd��4����3z�����I��O���GB�@�pFH�3k+�(�b���ẅ́ ��+���C�.�M��L]k��(^�D$�Io���bb�����g�~_?(�|�'�9&�_1t�6IW������MV����|���8���������� �ͮy
���������3|!J��Tg�:q��ܡ�!�i�����f�p0#il�ޮ��@��l1�iA,�N���q2E"�P|�>qI��O���2�kK�%�%b%������	����刈 ���G9���=!@�#�� 0'���m�>�)'��@���(�)N:,�S�"�R�z�F<)���+h(H�������Q���LȭZ>t�p� �G��&���m%��h�t�������\bj���0��j�E��
:KVq�>p:�
Y���	{�T�S1i���F%��'�13t�k��2��ᇒJo�w^�<��L��_���B�]7���&,"j=��pjT����٘f�PwLʷa�ĚN��k_6�\��`\�Ւ-�]���f;~72��?��޵��y�߻=\������3l�Lx�z��������g]k|��7�yZ��C�'�ͽ����a�
J��/���H��#]ݲiy��`���9�Y��H��{��i�LmLA趴��4��.s�P��������Be,�*kƺL�H�Pr��Uԁ���%1�ü��5���_�����(-6ս6���5��YVm�2���p@��{�i��N���3���]�>6�4�: �GϾ���r���#��������J��ᡷ91�Ѹ��1(n�:�?��S�~ۯmnl������c|~H{N��֣�3�M���/��wws�_�&[�@۹a����WGj�#�J���* ���]������
��Q�
���d�$��E����x���AE:�ݻ�*��X����-�L-{��̾hkb����;�-�a7D��'�����O5����m��iut�p�*�� ����,���u��&P�9�i�Ɋg�w\�uB�(�����b� gY�N����w�e�n�$�Q�Ӎt����{���3ӯ⥷F3��zk���rS֗ٛ���VnLTw4��w��?�ﺸ���W�+��}j�ӷ%:|��x
��G��f��W������g��ҔӅ�/U��1�v��*uI��׵��i�&��C��4�5��{��!L��J��?!��q�k�o�s��';��1I�!����7�2_����i[�cC�;t�I_�5��D�b��<��#��`�sHX.�aʪ�)�E{����C����ßݍ萭�0�k�2
������ע�����K������HsQ�t `�'!d�r7r��������d_���cG�����o��E�!��c2�W���ܷ���\|5s���g���$�x���{ֆH#.���)�ܒYh���q����%b'E��'�����h�(���@�* ,t9gZ����&�ځ��5��F�:�+�r��$�3��T,�s�2ue0�E�������M���=K⋆�=ܬ*��waCԘ��W�/*&k��4���~{��6xy/*���vҘ�S$>揟�V��~K,w�{�L�z���3�TͲ���R^V鴻6h���Ǔ>t�Z<���*B���2���3(2�Ǭ�r�GG���a�0�wp�˜ޠ���l�bA��=�ˋ����+�n��p����o�m.Hlr앜9��<ʛ��[y�`�[�> ���'Ķg,R��1��/
�����.o��G �Do\]wu0@-�/��w���T����[�/��\��k!&��3f�L��{ъl�D�������K��q�1Gj@F�p��c�ٞnȟ��!5��m ����.� �^3�닿��z�L�Q{���'cE�^���z��9�˻�&�ׂ�4�R8���7f��m�4})�
S�҈J�L��}-��3�S�&�E�ڈ�e��{?��@7�P�#��F�MV����|���u�x�䫃m~����,����.HE����k!y;Cg����ᶯ���i0��z�<��̯�߬s��iyO�c�t�@��G6%e����ۙ�|������k��� �c$å�G@ٛ�I��]��m��*g��&�g�T1��n��&�ɦ��&xa〝P�9�C��q�l�:�	�y�@{��`�q��@�-��������"�;TM���>@���
�n@��V��:���C��K/�;���i��m���ՙ�H�����^:M����H"��Au�-.�M^���[��X*��LL$�j�]8�e�H�M|�����F����C�϶��@ax8�ٶex�ˇT�$�,#�Ν��W{���iy3#�_�
�;-^;�`�Z�J
}CQ�q��6cd~s�m�R�n`��h�b��}���v���l�Oq�(V�s��/�!f�	����ϼQJv� ��nK	�|,��RMK����B�u�)���F��������xs����I�8_Q��*kj�?��K��������:�9?wy�S�8}����	Y��	��lS>M���sE�Ѭ����R{���`:ۓ����X��~��X#xX[E9��PA��x�v�H�t#-��s�� ,�x��&�


	YY�P���[����[��iw�(���}�H��%O9x��s����U� ��9Z����
�_;%"ϼw��!Ƃ�=��:�Y�L,t�F=[r5��g��֡��F�D�HAv&c4Y5JwG�i/��C��f�1Ǹ߂� �Ž$j��<�т9:�*�J�V��-�6>�lpD�[��-Q7Q���u-`?�9�1�Z���"�k#�/���ҍ֊�T4���F[�f�"�[fa��纹M�����C��e@�o&���n�;��H�QF���Xy�F���Z�oq<>�o�dd<Q/d,	KC�t\$� B�q'�KM�|�{�YK�ǁnt���ʸ� /${�6�"�[Ћ]L�_��=(��HSA���FG ʞ�vd}@��ԋ~]R)��Ҁ4���HO����$S�`]w>�W�h���4����'�����K�����;)Һ��`+s|�\��:�C;�~o1�����a�8-��	�$
*��Bgiox4��q�f��k����v��"!)7p:�뿳.ct0��̯G�Ξ��SMm���B���SB�#���^��!dk���J��V����������Tyu���q�)��J��`����9x����V�Fֿ����Uq��XW7#8gm�MNVk䜯n��<ۓ��Q��*滋L�k����0V�@�]͉AX�1 fUB������y\
� �d� �%ᘏ)"�͙.�G��OMv��C��|�3XUU_�a��s����$_��1drBxBH�nC��yI�'|'D�͹!��k���W E��YI�"�Mv���e��MQ'��[��Q)0*M�o:�\���"�{^ڊ��D�nҵ�{l�z���<9<�=��Q�����KRr|kG���;OJ��^�f����M��:�`ߩ�p\�04�<;#F&F����Cj����6�E�I�\3Lk9�^M��-��n���߭Ohq�Q��b!6BR�h��^�m'9̥�ݶ�(&gKb�c�T|��X;�\^��%����1�{�46u�Qe�K�ڃ�L+�0&�M}}=u�r�쒵ŕ���C��h�����}-8Jm�GksLN�b⥾=�56�ɂ��n�U�Pv0IC](rhz�����\Q/�p�g���͐����7��㏫�!��OG��Ф�j;*j��z|�r>���D��>1�C��(������bb4&
���I@�!�\%�M�Hb^Os��,����g?Q 6j�/@�cB�N"`����%� j�3��(�}�n/��k�?��H���S�%��\u�j��Z���$!ȯi��m�'=����p�� �j]\�;ެ����VRifP��=���M�1��������/�E�R�d�j�3�)�ô7���t�N�~ݣ�����-�~Qt^�Z��Q8���[�%�3�Qx��C����2H������x#;3�Vк1
5X� L!6���=�Q��Փ�U�N�H�O�M����]zd3 ��Zx��(�A��9����a
�ß��>�4�d%���b��`еC�L	n��	��e�݋Ï_1��A�dx��Ҋ�����yw�>1GѶ]�e�D|&�����a4�Kzbg���^.��b��@�ΤϹ����].�08�xhi�����I>�dF}��bm����!�H���J��"�d���Z�
�$�.�A�FG���"̀f_�הQ�#���Yjd�c��aR!"�hx���)yk�̢Mx�}��i띶��@�<�CB�@!#��Gq';E�Ȏ�{=��`Ad�#��r����yp�Q���R�NZ]b�^�>YQQ�#[C
��IMh'v}��P�4v���.��Oqz\�&Q<�{A?��e��A�����f��pdj����+(��ﴇ�gq�l{�7D\��H��-�Y>��){���z �&F�y�����MM�����">1qc�D�����ǘQ\Q_�6:��?�JЮ*��X�1��)�tw�ܺ�alɇ|�- �-�<̍1u� �羢�2����������v�!`4PV4�$B�P���#En�+����vJ*v_Ё�W"r&sLV��-9������g�`�]���5�.�/,��:J�PyZ�e�m*�m�@M	��4�*%�R��0��.�zP�X��^)���Fq<3ځ��L��_�R{���\�G9�U�h�3>�=��?̾B��)
q0M���hik�8H%*lU�����X�)�׵5M8f }6�&[�#�(��xʾi�~��R6�s�߹�!��p��G�傏QپlALx�6+@�P��+�J2�(Q2.^�����-�A\���عɋ&}g���HL5/��a���W��ڇ�\4M�V�CU�����s-�蓣[���Fr�����kJj�0U��&�g b<\��TCY}������w�K(�
;l�4�b��:����m��1f���}m�0�Hˏ�p�#�}��R����>�{{,f�w$��*ˠ
nv��,�fW���i��4���;�ƛZK�@��W�о��RTis��� ���փ���������k����8�I�4�sJc������Kȶ6�36�Җ&)���R�;���R8��~�����fr\
>�V�^�U"	Ņ�f�B���ﲀ��_Y܈���fE��z?]A�hOm|��Dou��'Y��4��u�ukC��v���r��2�/��f	��#����W�Ν�o^�F����|�i4]?�@)���Ɋ��d[��jdf���]�����"�p����/��[��7�����D��`�x�B:���m6��"׌���#�ч��Sz��yXe§T��7$����Q�v��d\�]������x��6���K\�6�aӊ��4ջg@���B�{��V(��	K�u�kHچu�nz������C�_rJp0>M,�Q0A��6o1�#$քe��虡3��^��#���I��޶�Mn˛_�oB�lCк䩁�˛:q��A��ՏG�z�$K�>8c�F9?+�!��)���%����IZ���
59q}��������p̮5r���^���ٝ���2��~W�qm�X���~~"�$+��?l�RF)Y3�����FR�(N�fx�*�����9"�\"˺�*�9�2�+[QU���WyI���J�Zy���1�z5�j(�7�J.l'��^ �����%3�&�@�Pxs��R�*�	���_����:�եR9�k'���cF�ο�涼g�{8}s��R�&}|�օ��l%��,y�.g��!{���B�Y�m�I��bA=�בaވ��3�im��ؖ�#�K��"����^��p`�,K=|^�`iYwdʂ&̼G��ń*5я��|-��R�l�f�[ƛ�â��e�9HMBe��#���3��_&:~<}��S껫�����Q��Ǘe�aN��L�L��m4�b%�1�8���{25f�]�35��.]��㺪���T�jJ��3��$�4, *��1�Ϳ��\��GD��_�����n�ܬ��׭���o?�g=I7�P~�� T8�Muo�?0�V �j9�n�&�%/q�����w�V�k��eν��=m�[̷c(8(���볏��'����B�b�LWw�+e_r�M�k�l����i<jɘ�دA R�z��8�¢6<¾Jt�z��4b&�=������}Z�^��N����A�,�{��(X�1��ddr��޽-o�(��D~���ځj���uC���?��jn�>d�k���).���}Suo�п�'��x���L	+�t�o��P�[�;O��&󨈽�o6���<BLN`�vwLY������
��=$\;�����_�o{��b.=��tLG�h��l�)��P�/;��TK�����M��`9���_t72m����L��gW�@�g�H�bj�:o]�k���� �⃩�b!|8�}��ΕJ��h0�:�٨xET���Av��'�Θ�g�ֳ�)�
�u��a�e�߱M ��#��I�֐�`���V�N� �4X`������?���*�MҬ�~P�H~(�5RvGKC��R�H�+�z��� M��Sbٗ�L��x�4Y �7!�}bEƐA�~B�F���T��UJ�1挶��xK�k���c�m�	��J��X]����OI��L�nUD��BP���7�{;S�.[�Bh�>`I�*s8r��#RvP��-2	�&}l }3I������q���5�>��3�l�����,[*�t�*u��W��iVoT������m�R S�8`j���"���ެ��^QiW�Cn��� �,�\p����F�kV�s��8��=�p�?PI�p��Gz����5�h���E��I�U�C�^��yt��%�B}�����lz�xrD�j���'*�ϒ;�?�41�:��$�
_X	�tc�wiHV\|)i��0����K��礒9�Gv]��tk���'�7E`���}��yZ=�U=�r�]�0ҡ��/��?��}�V��e�)�H弡�۸��l�����J��i:L�}����B���1�5���}��=��To�@�}*����pJ���7��Yw3v�;6o:X��5k�'�T�c�:uIk��QH����0�*�
zr��&;$FV���T��n�0��s=���7o�P��z��C='�U{⌧R=*@��:\����9�Q>��� -�J�h��z̄���_$`W������9�\O�bB��z��<LdB��q��I�g5�'�]�t9�'�T}iM��87�e�ƶ�H^��Jx�A(�H��F��-Z�K�Z6U\��Y���%�U'<���{�����+A"�X�N���D�~��y1f�q��f�g�ThW���Ԕ�(�&�w�v(E���w8�5?����2,Y�K^��p����M�q��UXt�֚&��/���.@�p$�,8W�*)��e���%�]�âQ�ͻ�C�?��@6R�/�lo��۟�W��?n�\̆����Ř�9�ۖm�;�G��}�R�����`� ��jz������"���N�'|�ؠ�W�b��)Uu���h���
��t=�tt&H��φG��Z$50��+*ɎH�Ӯ�Z*Q\�Ax0���%�y�>6��~� Jh��8��O3w`�[�uL[�K&g��W���CM S���<�
1�߼���0�a]5;�w���˧�0�d�ɇE�������F�i�}��"q>���O�SdvZ7�?�3���MG���}(������>*}�ς��	?��[�c[k�YY�	�\�6]��5"���f݀&�GwE���Ǣ�ې��%j��g�4h��H,��tG�ĭed���<7랎c��������;�n�wP|K�/.:r2�/����P����;��J�����#� ������{�('��H?C�~��L�%�:C�j��0~�\������E'������/�V� ��\Z1� ���4}�R���#��Inf#J{������6���|O�}]?��:��h�y�=�;z����z��ʏ��^�#/5�&��;\<WC3^݈�	�2i��>�P�~rW�I�"KI���M�T�4�V6߸S_<�ʋ�57�6�:��K8�'%�m}e>��:O�fӋe�bb%�u�9+V4w�H�~X���P��ܼ˿�54ts��]�M�2m���VHE�e..q�{���7y���BzN�����X�\磶�B�,+$�!*�<K��4�j�+�:[��!���s�PJMVׯӹ���V~cs�����@t�o�o���\B��nB��6&B�$�]��������p%4�ʝ+�J��U�R���t�̫�[��6�'=n��2�ՍmO�-����屔�혤��5�������)�c�s���]�S�Y@ʺg=�X�R�S��,wm7Y���\z�~$-�PGQn�=^��7я�#u>P����ظX��.�����rN~90c��"�����v��}�ƟK9+�0575Z�g⸡���dJC9�J�7��^ ɱ�>�.=�[Ф��)fp�o���v�?d��-2�}Q��S��gWi�� ������=����o�YD��?J�����{�<�U?��c�̙֭[�_hk�i�{�9�g��>�9!�	Ec'�c�3~��f�@�@R� s�C���F�QU�մ���и=J)��6����k��9I',kE2w����nS[�ʳЏ�J�zݑ�k��4�A�6��DY��T���������1����Zk���R�x��e�����7���n�v�Ms��0I�t�vkӆ�tF�Z�1EP�ż��pb*>PO;�ߕ���zdw�?'6�!\4yV�S��M���s��i7ӭJu��Y�.��{z�mn��2�ؼ��ˁp�A���ۣj67yb��>��\�� ��{3P������;���:�0ϡ�-�Ƙj�X�\Y��/��+���cV��0V���+.KA���C�x����2��T�����N�F����$�d��%��LRܘX��TJ��L�~���/�����G�*Ί
D�m���E�vβ��3:|�;}�~C�ɱ�����Iw��A<�%�F �=��)�`?�=Z�|��y|��$ 16Z��X=���)�gg����')0q�D��+�h�M�@OKs�3'����-$ �����(q}�ӋaSFac�[���e-!S��=����� آB���
���I�3lT5��5���H��FO/Ǚۚ,l�^�>�u�+(O�C�K���龅��)	oC���S���3�ڃ_z���Ư�{��/9RPӾZ���Wb7�8g.spO�eG�D���uu�Ve�>Q��VSͳ�����}$��6��.1�i&/�dw���]X����%e+������)��W�
��|6/�F� �f�Rd�n�A�;X��[�V-�ɀA����
:�f"3������T��>��U5���f�D�2`&��=18j�rҐ������C���u�������>T�}�����.!���.@\��\t�xQQ����ds���˯43$���K�C�|�r"4��e?�f4#�O}7E��W�O*cs�����$���M��k�O���Vr5�͖��[�=
�=\Vɺn�(�)H��u�ۨ+l�j.�d�&)��n�xf���AV�U�y�`צ;C^o�#b흥�2^�ň.��LFs��F�k?�n��J_��yM���v�'�~�3��e%�G���Z��m��U�� kQ�s���}M��<�?[�v_�����7���$��8N�K:ChY�-�M��3�l���+y�*;.%C�����?���m�߿��e�VePR���0K�h�)�(�e�(��B��+��k4�	�Jh�h%�-�Xn�튽��]<��p�3����罆�'9YAh��xgO�j��f�u�n�%�Y�]4��c{XӺ�2%���=Nո���T.m�%��2��9>Z���c��.�FcW�����~���y	Zt;}���i��z�:���n��˱H>[�ROǏ���]�9�r�d�7"9�4B�z����s+f�����IPYl����F��2&xM��$�I[Ǌ��W̊��i������A�Œ&�-�5iQ����Zq)j� =���.����;U8��m�Uv��C<eI\����C$b+t$���G�SS�<6]\�&����l~7a)Vf�6���χ*H��[���`��q���d��ҚY(.�IlD�9�v�,�v8��FT���#&���4�v���'��:���jh�(�NZ��uߡu����~��D�2=b����4ɴ�Җ�M����o�As���������/.����jL�&����������V�:��P��	]�T6ڪ^?c�Ӝ��nt���ݭOЏ�� 9�����nYohȧ%)�#*��%O���(NE/]̎��n�H��Pf�'�*h�S;͋�����L
��նE�`�uIb��� NhC��(�῝��F�֌)�+ӯZ�u@�h�aI)̽$���/��z�����c@>�c���x���@����o��,煴"چgC^x(
_�?�k�靽���^P�Z�(ΓG��ذ0��ȑ�W�����h�İ Їe��A�䣊��߬ѭ(��9�-�vb�~F�6�� \	�ƴ��ܷɄ�N�v=b�0P ��M�x��ܡsQu��c�tюF��ߗ �����d���K�&����D��Vx�	�c�s�۝ +��Ev_4�����%�mܑ�O��l����q�H��Ѿ���ߖ��"�j��-������������S�E]6� ����`�Z���f�(
a)�~���*y�J�ksY�\s��g��1���B�8ǟ�HvJ%ʭ���ȵ޿�b,��i3NL�O���1,��-����)By��+ٳ���$Q�p���bx��=�r��ս��!ʛ�0��[:ś���F�v%��P��dEU�>6�fk��zx$���e8>���v�:
h�
�)Y�x�F��wl��
`��%(�U���h�{ѥT�2�[@�0:q�)Ix�~>�Q�cO�ϊ��|��`�.Bj�
��~%UM)b�-�.��h��ա㉙`�2ִj�dnl*D%*�P�$I1�-�
�D�V�Tqg�uQ�~dU#Zy/%����M��T)�aI,�4n9yj/�$�G���s����x
M-���h�~��:*)��������ї���<��ŐEQ�Rm����$^����ʵaF���_�i�L�L�!rh5=��vke)��Z��c�5�M�^���.k$���J���� ���S�	(X����g��ٕ��b�\@�߅��C�j�G�;;e>���SQ;�xI��
u	X�G�}���RN2��.����sFZ	�f=��9#O	��REۗ+p�1�6��D���G}�2T�6NQ�<�J |���\�&���c]�Y0D!3����N��f��ڵ��y���B��K�쒑�e��ː��v����u�	<��ȭ1��/ � �956�[��ٌ��\��?0�80N�����c��J��v����t�#T'�DU>S�$џ��D�K�>����S�sE�o����eA���](�H�ٜ����2/�+��r��Σ�����r����~�C�E��I܇l��i�YV�F�d6��q��
�E}�f
q��Z#�a�����'�c��u�n뽝@L�WЗ�	�ZJVXe���6-�k���"���ߘ!�_��O:X�`�u���g��\\�e�
�cD�S|m�ܓ��ve�SEܮ�}*�$Z#b�E�7)-
���k�zE�ݠ�P��O��5�Ôuʁ�*��t�7�y��C#�	e:�Q����Z����'G-(GP�f�;��)3AA�H'n�>��}�V��سCQ@�QK8��*��{�! 򘹚Y��b�f�c��eRR\UA}4��g�.�7<t���N�w�uL��n���4(��0-����M�r�,���u���x5H���k&�
���@�g'��Rxm��=��"]��~�A^c��Q��>�@֖�q�vr)<��Yi�ih���9#H�y��b!j�]b#e0_�w��9"�Rhu����U��r���^�}e�,0��R;�Q��@���`�E�kȂVv�{�ZIF΄��?)sgE��=��S��W�s��~��}dxh_~Qk��PB�Cmj�#-��ոJ��"�<w�/�'|鲚Bɹ>����tcwb��V���hB^D*�\~�����pi� L���y� ��/���?��������A��>�ѕ@_�w&�	���׌�����H�'z0 R��|=O��z������ʽ2`��.�#w.�-��pH��Z.��u�3���pi�*fk=q�羽�W1ZnCM����M˪��eJ7�?�)sy���>�� �p9d؋
s�����T�g��V/���j_�By�_��!����q3�/��-��0>L��`bJbQ�F�y;���{�σ�m�&i��&���d�{�*Ɍ4�q�hW�ǅb�f��$ruz�]��''Q��pU���ڔ-�D����,D%�x�����G���W�.�u��v�%��cEM��I��݉��Te����F�}���T�HzI���d���֫�~�X�Cț���b��D=�1�T��|H(�����IT_�P�Y�ů��[�k��rY����a�,$�Aל��O�j��?�]�B���^�Gaq^�Ic��)'�v\U00�c�9�]��*\+�9��VE��F�$�*����Dv����L���e�Wg�7�]~Z����{���ep��`�Ո��l���N��>�܇��}^�����!q ��IqA��d�8������B�j�̈ c/f3OW�i�,�d��"�4�4v+ zUz?��J�oZ-��CF�ͻ����gcQC��#z�<�t�{V/t�r�� ��V�h� ?�[gB���A�fbO�rD%~���:�f �6�����	��-���Ex�ik�4�'��U��t�7
*0S��n�����M���ڞZ����t���&�ĸ��Or��+��{�Ct�5���-��l��>��w�-=��:�E�ס���ja��D�����/��{�J�Q��t�X�o�gix�,o׈��hs�!&<?�y�3u�����ɒS�f�'�"#b�7�.��:~Gqu�i��K����+E��2�@��_�-�(X�u*���9�aT��E(���{9K��_p_�������7��A�K���".J}l����i$٩(�!x]ѳř�K��$�i��. s4�����'I����MD�Wf�X_�H5dfi��j�˹��7�@q~1�i�j@5�۽���ןO ���Y��3\��>�؎�$'��r'�K���R"{���Ze8}Ֆ��oʙe"��S��+e����0���v-��g޻`-�aGtP⚽�cE�6)����S**�\�~�!V) ��;Sc�F ����k {o�vD�~�E���־�=/�C�æ�jlc0��}��#o��/��ħ���ٜ"�_��(�q��}0r��ܾ�ר�3��q��\��l�K�,F�u\Ր�w}�peM_���!��,mN�)�.���1P?؈�OS1�5.]}�?�M`a#&&J���b�����;Y�4ǅ���ʆ�����K+g�I�0v��G����{��̵0����ز�����P��n�� FX�{ƻ2�<��R����Ol%��N�~�׸��)�&yJ�<*�J?h-�@Ϧ��\5�~]��X��<I}�vq�\��޶�{�ǦtT�W���w��`cV�����8�&~Vu����>5#U�Ӈ����)y?4*
���˾t��9�dz%�㴯�	U,�gf
%�N#��Г#5���C,3`s]ƪ�x0-���,U��������W�uZiK�*�j� U�׊?3w��l��?��㣲��i����To��
�؍�z\��P�ȩ�P�u��)�ބa�`=&dN�OT�.h�� gV����`*I��yծ~��U�r�
���Љ\O����5���v�+��7o�
��4��m:E-����uEH���A��T�i�,j�Hh��1��t��`ƍ�Iw��QW��\�������I�_���>�ce�9�abK?�s�В�I��Ƹ&�Ϩ=s���[)>�Q
[�G�z�@&!��v����ٟRy��v�{��/ՠT�2���k����U�UW�qWj��XH�5r9�Yl�R3��� ���-ي��Sn;�^�0Az�P���{�t��p��c�v��o�J�^�g�$b�3B�a8J��R9cU�P!��ƾz�,:}q&��D��\4w3����g1�^�h�#���6i�_���g���@O�lG(�lD!��ct����aP�9�:�c)W"!�:c8�S��Ti����$�$�����uK�2�8�u���� ��,�-����wz�(�pl�ӧhuSN�8��H��Vā�$�ne�P����ӭ%�6}z���75B�33Sl些nh���Ӵ��&�$d�����:���Rj�V�l�[�N�e��+���q�����*�����5;�Ǯd!�tx}��)5�Ҁp bo�hZ��)���8i�`L��u)�.R �Lx�*8��/���j���g����&���h4hꎀ�,~כ�C���R�^�:��COZ(��1hB�bV
(�Ag�!�u�<�@H�պ�d�����ggK\\,��+��۾�;�\�p���P5�'V`SJ�Pv��JC�BX� )P�I��잌�p2��yJ��RF���u�ϣ�5W*"���lN�۞�N��C�7�Vx
�vu�"�������'��s;�3?��=g~�t�x��U�A�Y\ht.T㞨�:���u�@@�(�p�py�B�q5g2��{`�\�k-�,��3߁0�G��t	h]`2Q�RsJ�9���!�M��SfP*��hj���&T���Й��*l���z�% �y����0 �����!�9��T�V{OW\s$����*�O
G�()V�'��e���K��5��J� ��X.�<���I9�� ��F�K ��>�΂�%r6^�ʑM��~�}I�!T�}AzN)3(i��u�Kq�`����Ҷ~�'��Q1k��i�H6��G(��=���PvsK�i1��!��nB^�a�[(ÿ�`���w��ZE!0��0�-�g�΁|���������Ρ,��Rb2��9"!�<ˠ�L.r�����+ABB
���[tmkʲDYpΆ+hc�`�cQ75 ���5��[m�\��w}�>ֹm����>O��L���KΜ��P(��}?�^�� b�E~�gu>���psb���a�+Y1.����IBix�h�W~�D�c:�a>;B�X-kxgq��w����Ç�ޢ,g��% <�30����nc:-�!����^ū��
"c��P�EH� k;��+�uZ�5���J��!k�Z-qzz���G��Gu]�Y�	�    IDATm�!���.��OhN�����WE(>�P�OLF��A�"�UxĠ��B6b�-�sp>0���:��l�<C��4WJVy�,�N�X̏ص-_@)�</��Ǥ����S������r"�|�  �e9�"��\0�)r�P!�a����Rd���\\\u,K������S���.�]7B���A ���CA���JZ�6zN{������-���0$�F)C���
E^�(�������R��h;n�*�y����Y�Ag�ʠdx�<+1�.�e9���z]�����Q�k���u o��DY��^�X���eY�Z�����,�L����D�l6CY��JaR������:CQ�(��5�a��\a��Q���'Xǀ"c�=�_Nt�c���%�	S������B��͏PH���9ỐRB*��(0�0��h��B��pΣ�: �D�kt���-��)&�)@΅aa��:%c.�K����X,��=���B��B
��B�yB]��{#C�th�G0ƢiL�}j�i6�f�
�#�m��#v��{��A�p/�:T��[��;�P��O�IS�MؾQ��dR�>s�pl|����1�4���l6OsL���Y��Zݶ ��t
�%��UU#/&�Y������
�R N\�j8�qv~�z]�3]gЙ�i�$�3.��m����`�Rx�������W?�~۷��o��|YV��;/"�K��AU5a���tZb2-ж��F���y��5h[��3�D̋YТ(��D�7��ʻ��b{�" �%�J��iЃ��=%E����l��ﺊqՆ���@YNz� >�(BZX�Nk&=���!CZ��9��9�ﰮjtw�B��k���[�4u0�N�{��3��B�iZ�����?��t��Xܻw��-�p�.�,C׶L�6-�s�6��UU�ѣ��2�^��>����@�tO+�����֌�}��>����?"�}��w��m�#�%�����`ÕO(����s������y#@K�qxTg:���t��zv�:v�j�γe��X�V�%���@K���Z�0���r	�W^���|�G��Gx�;x��;���%�	e>Ť, @��"����V �ᭁ5�(h��!<��B�uP�6�O�\��n���C�+�f�fS4M�����θ4b�ZC����x��������U�֐���>��?��3��_�'%Fa�sLyD�Wlz�*&@��$|��Cҹ�N�3���9n���=d{b4U���C3��@��_8�K/��������s��iPkZ� f y��Ag�;dZ�[��j��Z�tLנ�j�NØ�T��%ڦ��w!���-���j�uu	c(-�SE�7��&��v���J[�8�\O���qf�D18`�t���T�M��{#" R�� b�G�����h8}���r#/�7�E
��q�օ����{8Hd,3�f�u%ڮCӶl/ �u�s�ͺZ�@��Ai�Z��yƳ���e��ڦ�T
�Y���7P�x��u���u-��KH)P�ϑY2���
u]�v���?@S/A��w�7�����v�jc;�w<:�������֯Q7����ѣG�\���Rq���ܡ��F�!v*O�f��4�ܔrwζ�|Ta$�Y �)5x�s���z|;4Ê��o�Ď���?א A @i�i�1�.<9��'��l��9:7��(Т�yTy�J�H���"����mנ�+�,��ZӠ�+ky�d�uΣi*cPR����g�NfX,��a���!u������g�M��J�d1��.��R�f���'�����"�F�g&ͨ�X$ 3��чw�L d$�N����ȼ��?~�o>��Ǐh�������wB �'���R�2/����������������w�R �<�,y|��/���5�0?�����������������G�`_�u쿿�39A>BE³��X�A4�pG�?y��H����h��,�Ls]�������x��u�5���~r �z6�� �@�� �R�6��b����Y��z������=|p֠m�(���ŕ�t����-v�;xk���M���-8�e����1{�
 ,��bQ�޶!:���?n�aEg�7��H� �6S���Z�n��Tx~{��9�����2��0�!b�Ym�~T@�S
���a��驪�����\�x��l�9�\��!�Z����4[X�E�Z@���XZ��%(�e�����w�P����
���E�$B\�B!"FP���z��7H!�)�طU
IH�' U�W(/M+�y�1f6�G":�P������W�>�7�}h��sу�����7XӶ�6�I���.��-�1|�� 븲�΢7(�c`	P�%�p��*�Cx�F>� �pP0���q��ĵ NuG �Χ���O�	)<Dg���ÅX�c�߿��JZ��a�a�8�g��O�M@���e��tP�$,�b�#�1�h��)�އ_��G���-Odˏ<�&\��`��;<mף�:��c�+7��ϕ�7�C�3y/2�J��笷L��as �L�ɜ�{xbD2�"���|�Tr
����x	������+��5��8p��C�N�*��hۉ��8۾}���3Q�"й�`� D�4O�xo9��ة�0ČyPp b�W
<������ȃpA����Ӆ��9|�_�΄јt0�� !uTs
� �yoi��e�!�L��C���Mo੗����@b�U̼^����?r����?)K#nb�=���N�⼏��)�c@Hb	��OH@����P*���AD�$ݲb�s�J>'�glI@�0]��)����wƣ�D��|(��d�%�/�F=F���N�K �p^�,l�.����	�H�Bt�w�%��I�/2��b�B�(�⚺���Կ�Hf��걗Ũ���"D�\%���L��]�T�P�"�5�!�^�Бv��t���9�1q~(�WPѶ`¯� E>�y�Yz�]AE$f�Gr��3<���8)�y?��}>8��C� ! rvO�����%��A��T16#���c���Ba���)-P�q�,�ɍd��D�H|��ȹ=Ĝ?IE�.��}��L��C����$U���O&?O�D��dv�������|��!.2�\9�����&�L�R�);I�*Ӛ�(���j�dp�1�u�ٟ F��P��q�`Ҙ�w
�ļ0�*dn''�яc�t��~���CI���
E�x4����W�>��yI���ʡ��=p����nO:C$@S�$���*�ұ̮�I�B����7mZ�ύ�ͧy.�8�4	2����)�D������$r����{�@���v�ˬJ���������A+E�l\P:���w�`g�B�:�ŬX]Ċ!���J�ML.f��(1h�HE��HD�$�b�C�Kf1�- ��d����`q)G�iɴZ�p�7vRf���\��!Gv��_�0?��'�\?N|Je��Y��a�� �@���9!D��zӟPX?z1:�X	b<Q9xYb�$�W��PP�Ƹ)�c܆`[	 & �l���|��S/�Q.�G�s0Y���HS��E
	��X�G�7��.�ȩp����S����`i��C�/�iW}�����wy���O�|��bŉ5Fm�	��YÑ����H���ٯCK��i�4E���u>_�ܓG��>#IdGP�r��B�?o��ߑb5�g��DR��W�x����j�@���π��(X1�3E����T.�2@H�˨��J�nN���_d>��Zf<L��BBƅļ�GƶG+6y*tɩ��`E�ǥ�ڟ��*hh��V(���1=����;���`��@(���_���1��ر�o^)en?Cl�S{8�HD�8�M����,~D�'e�-�0%Ѡ�� =EM�?[cX<WH+uB��9"����`M�S��C�� �EUUX,���
EY�*KT�UŹ;ZE���h6��Y���{�.P�*V%��->~�>~��]��9;q����E�6���ɸ��>ӥ�{Z�g�� ��L�~��1�H�(^�3�H-QU,�8ɉ�Hŧ��]׃B�*�(��O����,�QB��BH���؍^p+���ZP�m��j�U��(Q�2�"���Q�`����
e����G���Rp��\.�^-�Eoz����:H�?��� rg��S�����[�b���	��4h0!�#�#�ƭ��{�;����SkꃊBGL<l�sq/JO&@��y��;#���{Ԟ+�oۂO��f�0�Z���6��o�
m�a�t��
��$�����3<��������b����Y�v��B�FUV<~N���Q�5
�s%�u!��0��f>eY��j�v{lw;�e������\y�������Z�  �,�s�n���n��e�L��
�e���	��;�Q0I���$���xEq����4�u#)2#�P�'8�GCr UUMcL3H�A�%����&a¡P{�P��н������z�5��ʲ�.Kh�C ��r���@Ht%[�-5ʪ�w�YÕC]-P��"9[U5ʢ�.[�Z8�QU,K�Pu��r%��Fk���]k@A�TUt�5�9?���4������aOv�'8��%��	I�cv~c�#����`����2��y���I�;���cW����c��?C���?��m�[㩮H|��y�P^�B�$�$n5�EQ�(kU��xT�CYTP�d���p�w��VC���`��d�@���b��H�5(=[:���=�؟T�o|�
��-��:�=�u��A�D�l�䬏	�[��t'0�E������h�R������f���Z�/y)<R���x\%��ғ%��7#����̡�3�|�0�XG� a�(�p�<)
R��ΟA P��I�!����=�1��!� "�OS�9;��E��	�z�]����}o@���RHD{!+9,�Eq��[��=��ND�s����?�Z�Ѵn>_�'n]��
X��Z��7�y"�����fl_��AuB���4,}�XB��7�Z���7π��z ���n�]�@<)1�E��s�B�Y���w�=�y�%$Ow$�o�o�6{�U�E]ø�.��d���m!�{4m�����C߶����� ����s	6&�Yk୅ ��	���@�6���
i�����v��ŧ���q6���Y4�>{�?�_�����}($�����c���iQpl�8��[�Ρ��r��R6 M��������[����aߴ�ֲ`LJڒ@����UQ"����򪬡�B׶p���q�}�Fi,�+��@����"����9��}��k�$ʢ�-+h]�4J��^UV�5� 
(
��P����"���>��L$*)q�E'��o�!'µ���5��r��+��Gx�8�82��瞷y�2�G�ޟ�~�
�>y��؏U��Hq!P�<c]Q���(�"�v;CȿFJvA����4�]P`��c�� ���;��k�bM}�	�� (t��,�����P���
��.6[�7W�X]b�XCJ��b��b���a,G�:o �f׋�ec;4M!6������x\����R���R�x0�M�Ɩܚ&�~����I��z�F-�1P�S�7l�i�a$�]d$�?V1
�lRL2�Op�S�@��m���{8��F��� �,����ث$�]ס�Z�E��e�����:*l�u]��j��7�AU��[]WX,jӢi,�5V����~�v������-'b�ObP,쑖'M��9�O؃@M����|
f����8����-��-�vئ�:���ᜍ{<������th�w���O!_d��m�)xg�{��
���c�d `Ct�O������=�٣iy�k�+Xgpww��i���^�y�-�0��Ǐ���~��ڶ��q�C��6*g�!=�y�њ���p :�x�gx;+e_�PĜnI��`Lc
t]����:��h���,�w}׵1l�#x��[��="�11��� �F�u�J��l��$�'���@���Rr;�}����^9����~����>V%������O����h���PU%V���[lww̡��� ~^�`>�x�tG��<c��9�<S_�oY��� !�;8B@I��(Q��B�{�d��I��9�]�sL��������u!fܰ1W2�E��$�Xe�|�Q�*xs�PZ�2����sޏ�0fk{\\�8�^T��,�����P����ݱ��9���_��7yz�v�����E�*�B�R�O��M����1�Yrl��莹����	P��UrZS���xVu��2�
�bL�1-�kX����MH1�t%�Y�0�Q� ��(�
#�0Z�b�-�p8��Pt�'boX�NX��˻_p���nw��n!ʪ���kl.�x���� cZt}��k!�Z��u����P�K�=�����t���<�X��3^�g@�O�Ƚ����"G}�TH�@`'|�2�d�`9�D����x����e>%�I�A�(�JJ�ȝ��M��ꃗ�ج�'o͍����4,�NB	�8S'���
��
�v�႗Ja�X`�\BJ�w!x��&Kk_0���|&�cN�b���]m�}���oϫ��*���Z9p�#z�@}�?V���ᬅte�99�jX��=s�|4�N`�!$A*�	2:�Go�(�DQH�@�=se����k��(�BY*�Ɓ������N��[��H�\�hRl��R�,�����Z~gEo�wm��y6Z���~��i@�\� ���x���3�R��Y<������Z�|�?���T&�#	~���E��},yl|�P��22!�A2��3(��#���d�(8HA ɻ$F��M���_`��9�\�, ��{y�0UP)���#@d��s	R�f{��X�/��r�B<�t�@+�}�G�r�S������N���N�U'��
ET)�s(t��	G��=�j�X��ϧ���B9R?��F�������S�"�(�%�Z���m5J�΁�B:)��>U��e᜖��e��s]]V�u�I<!���,t�&M(���Ɂ1� ����xW��z,��zu�}s���k�}��[���q��ʊ�v߳�-���d�7�H��R������S������ê�,C
G����b�|�{��H~
@��1zB��U�ɮc�5�.�,FQ��vjD >�h�bX��؄�z8�!�DYj֟�2D4j"�s�D{p��P	��a�_�A*��A�PC�hQT��%�*�=P���`�$Ƞm��n�0�D� �Kn�1
��a��&�h9�`�>�ϩ��q�IΑp�I���S�FFJ��a2yc ���|m�$I*iWÔ�?�B+Ǐ�8�~&���=}u�����i���x� �������@ ���R�PZjx����kST��H�
8�7��<�q�&d��-�QH��<��Z@�8B>N�b���ʇ $�تR�ZWXTk���\�F���X�m[�-/-���)���`u��_���=��iB�o�a�*�@�4.�NO��|ra�ˌwyxo)�m�$�������c�cz��i��=t�
�8�d[��k��Ӈ#q��'J���$SjAL. 
����E���:t$�@�4���r��@��
)$��� O�ʅ͠y;9f@�x�GoVp�����
��sm�Q5O���d��)n�H���x�@ÀR@�
U��f}�ۻO���A ��c-Lo PE���B��p1��Bj�+xL�"��}�~"��X�ʌ{��.^	��!Wm�k=p�	kr�����J`H	�A�y�9�7x��K��$nL@�x"�����X9ǝ0��d�B�J�U�R��G��L�P�1n3���Z�[�*GkLϓ�q�?��Y�z�ަ�{��K'1�uP2@Q�3y�*��u`�Hy����=e6g}���>��zԵ���u]@H�����1(�    IDAT�R���E�uxi�����>4�{�m18���^E�	�$��_�2"�π�G^��B��Dh2�v��B�>��=L����"!�b+2�̦'~�tz F<�6z�$�cؠ�Dd�`w'czk}0�p�-��\]��
� 8���߲k����E�����t� ����ѯ�d�#AӸ҈�ڄ��h>�S��XRK�󏔆��"gɑ4'e�,���t�'�IMw�o���\"q+�j��>��K%�E��x�����EY ±��qh��&�c����|S���!bi���KErUU���l�d��=�,٤�m����ϟqww�l,�}Z+TU�j]�?[�qg��B����)�<6t�88�*Ƴ1�6f�S�G���*e*�k%]/c��1�:}f�o?x�=d;�P��� ��(b��T���n�(eYN.�|91b�͈e;(�p�K1�)I��.19U� ���"
PZ�,J,Tu!�s0}��c3���@ v���|�����0��T h�Q�u�r^V�3ڃ��N����+2Y�<~(Zc쁒�$�g�M�~@��_R���D��s��q���<tα�j�,�}V����'���vj �z�����5��IG���MA	l��� ���syv�-nooq{w�C��̉�I����d���I�e2��S�����2�1���6�O���埄�q�"3�"J�-��|���<�w<q����r����TqᏗ�fO�9ȱ�B��Z)h��r����(&���m�����ڮA���s�P��&���931;<���7�Q���&����s��^T9=�8���oԢ(��\��v��c���"�i��54T)B����2��Ǳ4��9SJe��(
�u��r��(���{�+(-G�
)8�����t��6W2���d�4�J'�Ñ�倛f�	M�z&�z��U����g��lFME��M�W0Ơ�{�`����W@��gR6蕎�;���Q�2m���WQRHP ��U��D��b����^�pyy�JHY`���oQT���_a�cXסm��u	!*��b� e!ً �(�AZȚ�q���-�L�-c?q�_oO.����پ�]���dD�M���R�,��'V)6����B�����0��8S�ՠ�3�(��3�"��[��b��f��j��r=dK$�?Gc,D�咽]ʘɜ��2�:UpRD�I?�8~a`r��2�F�ibơ I�iV��H<r���H�r̪`�#��U�Y)�"�&.o�(a��h�&;ߧ>�}Ԋ�OvBp����Z���S)H!���3\��5���߼���o���;\]^A)�;�R�k����-�m��}Ƈ�������s�<�bG8���	�d'ڕ㾮� �|��T)����9�X��9��ҟ��*O�`Wz�49��0��M�	��l�����8�>
�A�I�d� �]%OuV��}�޾�^�z��r��R$Y�7 ��M�ps�?�����g�v^$,�=��_\D�	����Ϲcۣ���~@9Y�� ���¨J~�t�����RY^�RB�Z�f����:�\\`�z=R)R7�8��ձI�$#��,�E��X)(���&��\]�ƛ׿������
J����� ,W��>���:�p����+���ӞZ���� @���Q�EG��2��2���<�3�x3�(/�,�Ke�[V�!O%JU���X�v���R��)F���o�%lB����J@�eQE�]��Z���5^���!��0�$�g�.@X�����Z���\�PJ�9��}�m���+�uޯ9mZ<�rx��Ϗj)���PB@�B*������7�Nj!PE�+��UU���&������:&��$�y�x��<H�ZvQ���l�^��Z��T���Wo�^_B����4X-��"n�J`���v�O�>`��Co��s�0��"8���张r���N��S�&��Rȃ]+�t��>v���>>����$�?�Gz�7)��y�� �{c!�1���1��KUJ=v]�u)ֺ�Hj�מ�L0�L�#~���VXX�%ɀ�X�py�
WWW���BYV(t���+�W� �|�n��P��Ux������/�m����Eބվ���37
�p�^ҡw����iM���Z��s�C���c�G�����-6~MKx[�u�x-SU�2_4�Z��{ z���z��b1��`)Z9�4U/��#�1񫤂�*/��,�/ (FzT5{��e�W�^�ի�ج7Xo6�W$5 ���-����7�C����n~��>~����M��в$��>���C�R��m���)$$?G�s�"�Q��w8B�G��9���d�l@����V�󽞔k�6�E�q3%��8йx�Ie����_�J��YX�P�5���4��y�/)%��u��B����t
! ���~�p�G�s�|#I� ���l�$E���c���������DUV���Kmt]�ۛk8砣J��Dww�������o�����٢�Ӳ~�
'�W<3��d&7���RCK5i!�Y,��;ŝ�(_Kv��N��c�����	���]����X5�1/�3N�nc-�d����ޱ�h�A(G@]��d�(߭��2�&�E3�U��F��R
��!��:XkQ���.Xk�w]oa��d���r��bOL7�Y[�5.��p���D,H"�R����Rj��k�U	�,�nn�q}�	�����ݡ�`✁.zɎ]־��;��4Hُ���n���	rE0��]���g��1����ɁcBtP�L\��*� �f��q >�zr�r�򼤆����Ǫ�L
�PDk��j���Kl6��������
��������������Ǐ��mwx��W���W8�<�f�H����x��6� `z�i�Q�5@ְ��իWP
��������n�>c��C�60��w6��8w�H[@_*O�zL��ӥ���S�dOƎF��R
�ˣ���|�Zk�^3H>���В��O0\8ʷ�O�>�� �ǏJ]�Y�&� ��{�F�bX$"\\\�ի�����z�W���d��� �Ļw�b� �D�K�y���}c,��X�7����1�88硤�Skڶ�~�D��Q`�r:����g|����v�;t�m��
B�ˈs�'��V�����S�c��~L�6��� �)�w ?��ִ"�?ǘ��p�E��rQa�C�ծ�����Q�J�l.��~dQ��rҘ/O|�r�(_T�y4�!���Ѻ����߿�R
��
Zi�~���
��"Z!��hۖ�z�ݮ�s�n-�*>X��a@��m���gծ�o|������?�mwh�=��a]� ��f��\��XM_�Z��Ñ	����?NU$�B�c�ɩ�Uʔ�q�E�����yl�rڝ�!o��(!Je�������}@� e�Wz�e���";x	��K,jV�2�Ig�aN�X8磹t3�K�@�p�ŝs�1��'R�q�M�E��Л�t�d9�P*J����� yo�c��ȍ~dN%��sy(�^����X�1����'?[ʃ��Y�8f�tL� A������/����!HC�!�{7L�,?��b�G�Zf{Ȯ��u�U��nZ��b��R��F֡����$��eU`�� Dh��:�%�+%PV�w[��-������amc{^�.���>�Tc=V�Oƃ�����}������8�J���q�%|���L�yړ�r�7�O�$�	!��5AvHR��Aj_RG*�B����G�wy�B��EQ��*�u-��@E�V����P�����z?���(K9/�]��{���1��g��t��L>�q
�Rj(M%p�I8����/&7���C�^��8(�F��{ %����i ��hx\�L�)%�g��<�y�Ŋ�L8��5�lB@$�,pSQY�?<�v���a�٠^q���R�z�@]�h�m�GU����X����
��7�a�ۣ�Z��N�׶�v�-���������(N�6��&�G�6���s����|�)��s��m+���p���=>������Jeb�nm�G��Z/�X���!(-�^/�X,���4M����������ȩ�4�-O��ޠ�Bm$9D�O��m��sUT�2b��H��R@)-^��ĥ3�<�ChX!���?1����� �\�|�42x4<v�JL}��0��@Â����E�������~��! �CH��(t�����vw���mZ4M;C[�`��5�lzno@L�'��bQ�>�,�<�H 
>z�<�s\������B��O��Ǵ:����omjm��bǬO91J~N��H �I�ov��s����F�Y�H���1v#�,eU�(4�R���zӣ,h] ����ۦ��۝�nk]�*��ϊ[gy q:\	��̬�
���&a<=�$D�_a@�g��m9�D�F����ڊ�\����y�����=c�3�|G 9��(a�[q��p���ӛ�q���qڢ;�մ�B��c��D��ӓ-x_��-��j^2q�� (h��L�Xk0X���n����ɡԠ�xګ�X�5��$��e�#��!���)�����������'�����g�9�ƒ�C�R�iI�(Ox���L����ୁ��Xc �� �Ja6�fae1o9'����,�V p"��e!QUU�m[k(����v-�*"�B�,h��
�܀in�D��;����͟4DiD3��?�� ���g��[��Pr���=�"kƉ I�L���O�����:�,D`��W�SY<N*m�����E~�=� <�OK�ZK����Q�碑�}z��/K��=<��>����"��ay����P�R0�P������8��fv����C������EJj��eG/�#ϟ�S������z��@�;�?�:ǚ�Q�3]kyS4��%�6.`�$�flDM�՝!z�$�#�q:���zc��+ԋ
E� d"���hxQW�(gy��'<ȏ7��bncy��e�#�+� �a�8���	�� ���Ҝh������O����8z����h]�?���.�K���[�g�I'&����F;��H@	!t6ݡq�`�-8�O1�!�x�q@2��m�H�Z��,�*
�xt�E	�4�ȋIVr=B@�(��57�d6|"�D��V<TĨ���dב��T?�����2.��$��x��"w\��H��W0a��̠�fm�)�1��㏪?�)8�$BSJ�πA�|I��@�r$��~0PR1�8�)! ��#IMZ�l� �b5px2re���WBJ���m��v&tI@H���qT�˜�(m�����D�yB�U�}Uɑ�������b%4ӌ���o�n0�M��4� �	*>gD���\i�7|x�8�Ĥ(�
B�h��Ͻ��	�W��9�`L���(��+&,H� �JyF�b���F�cN����f�׬����P�ɨGd%ݬ4�����~N� �.�!�@$!FI�D!DQ\H�!�����o+�͗��BL!������>�L��Z*�{B��F�9J#�9H(I����%!��4�����G��d�����q;�
�iM˳%�|�#g&���7��RP������q��6�� ��xB&���1/&&�өh;���8Y�
�X����(Rf�`0I�$Y�,%��$b� ��s��"�<J&zD�#��a�G���d����R�m��l?kJB@�M��s..�hE��,�B��w �Ie ��I� >�M�E�@]/���8�u�7�_C
�����3�� ����=o<���#8<�u�c�V������#��8��ʛ�:Z{�	!����,}!���ό$~·��}��c�)��b9M�aB1!~��!�*V�Z-���Z'Cm�Z��ʒ�ҕ�BA�eQ!¾i�\�cdvwӪ��wƿ��x���j�	���������G���Gd�l�zY�V`���Dx��~lR�޷��. ������V[����3xZРAQJBN���
?�C8!�nc9��Ҩ*��x�az�d�Q�
D"��}�!�d���RC
��(��@]ל2xy����a�Za�^�9��C�:n>��>D�AO�>��9���[�C����ӛ�G�Q��џ;��I��X�?V�N1n}f�%�e�In��(/���E*>M�z��r�����.�{�'?>�F������,�r��8�ԕ�6.�(P��X����{����������}�C²��t������E�@Y�x��=����R
��>}��FQX��~.�!���ǟ���O��-����t��Im�S����<�M�Y��%O���=1;�9Hk���w!J�ʃ��h x�1�ESq��I[�*�ʉ)�J���[ ��1>�(H#xI�J���e��r��X�5����o޼�#���7�	Y��&@��Y��#s>�t7�`-����d^��nuNW(�b �"3����(L��	X�s���0%NS
,�K�B��*�.v�[�xg�%�,��H�1>ၓ1B�09.�K�Ah{���\�Z���]g`�E�,겄,$J���e��r���K�{�'�{�.������*�f��g{ɮ�bhz+,�g�6<P}|��p(��F��t����4���>�3��w�- _��4'����6���l�X�zsp�:p�ǰt�A_ e�� ��h�s��n�Nx�3�$�=IY�P
�, Eg#!(J��WWW��\��+,K�y��_�FU���2�u�)�Dn��,G�	6oS��5|��s����Nc�|n9�M������o�+�c�t�g��"��:>[@��7)���������c�DU׸�� 얶�qѧ$�H�r�@�ӦS��񌻈��e�C �� �0��~ߢk-/J��Zb]�0ơo{�.�����������a?�Պm$���f���&�s��X,�Z�ж{�v{���v�p(_(Os*�ӛ�@�����1�Y<a��\�p
�SV(Cr e����Q �@%��%�d�Tƌ�ta��]���>g����o')8ldK;ъ����	>V#J �A,�RB�Z�����%..���������޽C��QvTS�Aa>��&:�q����+���rJ5qߓKOQ���O͔�'�X��}7������1��b.ٟJ�[?̅p��}A���E��1��Oȩ8��*,��r�@R�8g�Zr�b�"^
E�QO5
Q���-�,P�
Z=L\, U��wu��jy�w����������7X�X�P̇���1�����xK�Ph��?�Ǐ�c���{)꺆��x�ه@��������㑥��Ɓ�ǴIJ��5�8��h���r�$_���Ui��ּW/�uvJ��=��۳]�p�k!��Q�Ő3À��d"^B��^��w ����\�x�S�X,V��%��������5��=����J�h���1u]`�Z��z�v;�v\�䠰���<������1ϓ��8D�����%��$d�<�B�����gly����yʊ3�|�7�8m�*�E���S��3�`J+Te�b�Jm� ��e¼�2(�'8�%2Q
� �ِ�ƪ����o���;��z�W�����3�Zc���Vt�t��w����+�Yk��:H)���[(%������7'c;�2���J2\ѷ߶��`/qĢ`\�$ :E?�ss�P^�E��Z��U���(�b$f
�͉�z�5\����U�{}a��	�3�6����<�`�s3�PJ��j�y���_��������_���~��#�9�=�6kH%��6���C]���2_��Xg�Z-��훼�ֶm�A��<�~۟�&��i�AS;�*�cG==�����R�3������(/��q5<U'Ƙ��&�(q��H�^��P�*ж��q�=�)I�C����r�ƫW�qu�
�� ���ps�!\^n�%?���S��_�?����M���|��M��~��K�6�#������    IDAT��Ǹ^���� &�}O�xή�/���Q��w�O鞭�����s� �Z� l���c_
�XX�X�����9|���t�I)�U�������?��Xc�u>�|�j�΀�u})�Ţ@h�=>����oѶ���1����eYf��,5�R P�u2�
�룉7��3դ�G�x���g@��%t�i2-�����%����.�4bbU���FQ,PWZUX�/����ޢ�{(���R�H�
	�U
]@J��,b�HF:8g`;󛾝�"��[�50]�����g��e�[k�C.�ɀ.4�$�������G�������R9�3��R���Ԧ����v���_�7�q��_��O���K�Bs�5�L�I�<�2��L�3��|i�I�6&y���b>s(��h9�d�e��҂�E3Ơ7&g'�]h� E0P*�(
�*���z��ԛ�[K���7?�E�Vz��\�5.�^���:h�#	l�X��*����c6����kY�πb���h���Y�漍 B��FD� �@Y��G�<E{0�Û[<�`@	��^�4ԈH�1e@+-��x���}-��Zhcb��"��m�-󰦑vÊ"�'%&��|��=�� ��G��y�e&��J �P�Qg3b��B��;P6&��Q�;�$R.�V���ZUX�+�7kHQ��Ϻ�~�G۵�B���mE�f��z��r�@�X�,X_UU�7�R���!��.$������4;�m����u����Z�|�
A�L�\6� F7��6��9�����ϔ�xv�;!����10B|�d$Mt�6�z�Ov0�
v�>n����C9?�{Gń���	s��`t��﨔�W�xg� �($ ���%kE�5�*d�}��p�=��PR�>�sX������AJ	k��%޾}��,���p��r}��z��m�vmt�W(��%��-���1-W&=�8���tJ�<9��b7�� ���Y)%=V��P��<б��?+�%�Au�'�Y)���-��`��.H(��&[G!4����~t��f}g={fH��g����WW�"���iQ�|\�0���9c;���u=��ݣ�����1X�Y�&MUI�MԺ�����M�*V���z|��b��w��9L�T�%�-��/��J���#Ls���9,��0+��9�P���@��{�]��+�Q�kH��=��z� ��N�K���6��� ض-���z���PU,��t�1�z-B𸾶��nr��4;�v[�ɂ}o��[�]g}��dK�����9��� �����4���;VP��%	�t��ӛ�.�BY �@.<?���*]�J��L��B�j�E���X.L�ج:���;��AJ���lh�[��j�K6�.���M����GX�c�X�,KXg��M6?����C�2/c���> �J�����\h~���'��<᏾'��3W��>�C��HL��%U RJ� F¶cv
G�QoT����cYEg��˞ ͽKƮ�D�	ю@���[x'�t��)����ƙqk�\������}�}��,����no?�Ç��_�o߾�n����>}���'4m��ma��vl?��s6!�#�������%Y<\��{ ��T��w<� :%l��R���"Rv
"b�&7_Ys�<]u ma-���
��
}���� ��Ȉ/��7h����+޽{���O��EQ���Ι�;��~��-��0tcz���#��xo���rFAN��4n�d���0��y���>=T��?GG���Q�+�����N��8��<��y��
a�z���WL��)��1��������ߙq�q0�6tr��X�v�@Ij����*�y~�\BF�&���%�� ��Ǐ 
���  |����6������-���~��v{�����n��F~'#�\�hS8�f�!V3�}��(�dv�[�|�j{�����e�q[3�Y�{P���anr���tJ���tg�������ۦB(z��$a��~��Z���G�̛���D'���������.qyu�����o�!��f�j���`��������̀RUE����Ӄl\���d�|~{ P��;���/��?��P~,�9�"綈e�>�o^����/�h���=�Wu��z�����{��m��Ш��ָ����n�����-( �����a�g�/�z#;�����&�v� ?3�:V�$k��S��q���i%G�ű�_<�����$�{P���)f�l|O� � �������C��X6x�az����AUi�I� `�la�~�e��*�Z����nG����J�QU5t��>��7�7;tm��Ը���e>k���!��+(�F��Xk2�y�8[y�gr���<������K���ÿ?�|f&�
�W�s�d^��A���Cy1uk�G�r���}��.�5�E�4�./����<�87�(4������B���?��6���%�R�n��[����������v{�x��q�$Q�U~���D�xT:��ce<�f�&����5!�N���3�G	��^�f�} �-�pP�d���m��y�zJ8�������/;]� ʘ�su��%eY�(8Ck��, �@�l��o�������nooQ�L�cp}}!�w���o�+��?���'|��>|� ��	R*E"�jZ�s�`�-�O�����t��cH�,U
=����AmN��,k�pbB4��=�$p�>�K9�3�|�n��>���8���e�� J<�����WW�xuu�n�����RC	
Ig�<�.lI`�&�s��o���k�Xbs�@��}��j	)�zӣkۨ����FZ������&s��gk����f<
�#ؕN�)A#��t�ǩ
����;ܱ���ȘF��'-
�Op-����;���)󋟜���������Z=MXR}qq�ׯߠ���ѣi�KVK��4z�sʠ ���lvd���
��`���=@M�`���;��(�^����k\\l���+������?��}��ʇi�r.4��4t,�����Q�����=�.}�Ǟ������r	_���ڝ(Zk$�^���m"�s��}�d��i���pF�4z�R(]��
���pyy�YjϦ�im]�!��жm&�vwp:u�����I�m�@
UUa�ހx��~����@�P���O�cK����)�RF�S���K���ppZ�{���%�z'1;I�b~M(J�Hh��c�WT�-!F�C��a�B���t���G<��yK�{2S���e��f������#�F�=N��`�~ny�+_�$��(No��@���J X
��M&�EQ���׸���r�B]-p{w����E�7o�@���]Ѳ�@4䩪
UYfϕ�r�W�^a�X"�	*+�[�(t���`M�zu���?^��/�����;�Ӌ��5��$��(�5�ȒpEGc"61��_xIG*�M�DHa:�DS�A
�@"V�C;0�/d<�S���B��H���+�b]^���/yˊX��[^�����,
�V+���_6>wJ9H�Ps\�������N��I@�&�"!��68��v��d~Ç�e�2U&�����%�fs�ׯ�B딣��7�����5����n���1�mע�J�%J�P�>��K�u���v۠��� '늭��r�ƻ_�a�����-����w��P�v��O71�|��E�a�ʄ����`-+i�+���Y��P�D���+	(R�cY�Q� $EBN�<_H
�[ �BC*�]�ؤlhk]����x�B@�!����AK>p҂�"oT)h-#�;��(��J_��~�����1��ӑKU)9����M[�\�V@(�D�&Ԉ�m��ޮM����777h�-�h���[��G�6��goT&c�a�ƶmqw��r��r��xQpss�������+���^��:4�?~��O�#��E��@�����w>(b(;��	���������ς�1���Z/1���f9k�8�}jR�'����1)+GT|�3y|���lz~B@!x�rƱV*Jgzx���(%�Zk��	LD0�������EjM�9��7h�=��b	�J���O�M|&�׺^��]a�ۣ�j���Ϩ�E�����;t�G�e�7o������h��.��&4����7��=��*�f贌��(��G����c��;4�oHyIO�8C+cc2At�s6��<��#_��?����?���S�P�|�r�(ē%��QX�ָ���R
��\M4M�9��ni|�n�nq{{Ei=�Oe�p�;�`���cXk���l�X�6P��&��u��\B�>��޻������_�޼y��}��ϟ���oh�=�7�К�b�?�/X<T��o����l��E���Zg/�����:��A���O�ۙQ@QT(�����R��L�Y�ħ2|�Qq{���nw_h*޼��,��ֳ�(#���Ư^��f���\9i�2��5W*���Ko к�_������]�����;V+>x��8Mjp#�������c^�?�E�"P�AߤENN�y:�$��(�P�@v�s��g�����/���I`��Q$Ҙ�/���������7�rcI�E����B����̪z���?�/�K�����A��oSu�NeޅK, ���537w8�� � ��y��.�***r}��b����$냸�m6k<����m�^���NZ�;���Ke{:͔��;}����>}̼��7��o���w��Ck��r��R�l�TU�H;<FWh�p�w2�h+l�m�A��hy	hS>��T�Q�3(��Iz_�`H@�Fa�n�PxK��+$�e�Ln��;f'T{�I�P^A�"������P���g���p{{�E�ct��3�A��'�L�X���B��}�d�h�(n�:%�[rsKZ�$�g����z����t������Z�w�~�7Lx�D�v���B�H�յ=@"�Z,�x��-B�h6u�h�h��De[Uu���8�3�0^:�W��z�vn�/}OM'KPI��j,��-�Ez�J�H���E�qF�Օ�!-Whm�q��DG频��]tU��q��s��"��#�����i��B���8�P�bԂ�R����w�FG��B�n�}�b� �����a���r��`�Z-qw��h�^t'�����ݤS�Z�j�]����Ծ�����\r��O]WE�Ю��4s�
*�#�������������rෝ��t2��j������
��uS�(���{��U��u�.mam�?��O��R�ţ�@�z�8=2�ZE�m/�:S�H�Yk{#�u�`�\���>�>�Zhm�\�؎؊�m�vۡ�~B�,P�nn����-~��7���f�m���]�E��\�!C����<��pl"���e�_�R%`�E]Wh�zt~5�Fz�u������B�Z���&S��`�P�U��J��x�H��:#�Xt�n����:�9��&��s'&�@-O| o0*_��*V#m����=LU�25�z�M�e��Q9�3%.,��9�>a�lyo��{Hڝ؟��ZF���5gn��|bΫ�/"���9C�4>NUձ��S�����?`˃,�ֺ�	Y���t��m�	O۶�l�^?ƭᴉ,��N(ɿ��N�/���R����bH�Q�;f�}c�<��`��7Wop��F�vxxX���noo�����Ct�{@�mce#���������A+:��Yo�'�_P�@7�'� R�����8RN�ڳ�kF���?�ǧK���F:/��`�K;��ߒKk{l�����:�]Qx�p��	�r;P�G3����8% �6Кг���Y��0�����ĩ�`/���q��y�Օ8��}����?�����`*Y>\]�"��ܐD�#8��q@^��;{jv�������ce��cI��nP�u���Z�F���ڧ�ߏF��Ǟ��j��Ny��F��1�In0��&���b���6�ѯc���0ZC+]��V �l�I)���8pM"ƒֹ��s&/��#�|��v����͛[��\c�h�4�n��o�X6x��{(,~�@*`�}�%�����X}����2�
7�ځ�/�Q�J]׹}������2C�j�(�P��i�:��	��|a�̙�׏�;�Zxo���D��0�H�%C�)����G�q髮��΋(��8�NN�r":o�}@�{�>|��j�B�H)HKsu���7ר�
}����3�֑h�J�'���	g�˗��O�Yc#�E;�M���� m��׸i�e��*���W/x�.S��jI䬜,]�ɶ���Zt��9���H�@
�睐rY�W¥��|U�0*�d-�#!�9�ULn˼��b	Q0(e2wsw����
W�en�z��	~��w���w|��1>�iV?MJ�&�a��\�ob��[�w]wz������b�>_����~EMH��<<>
!'>��'Rk��
�9j!����CGe�I��,��6��+Seæ��x�G����]������ۛ[ܾ��j\��;�������?�z�0Q�����r���4��c�m�(;_�|�@�2�iR,')�$�D[Ҷ[�k� �׏q�2�,*�CFL�� �.�Dȉ .:�ј�+oȴ��Z$����V?�b� �4g�/DP������J��}��΢�[0��ڐbh�L$�^��J�CA�Iv�SK��|�|�4�KS6�i,h2ug�PN�7Xn9r��͹E�ʆ���8&�F\E��4+��̗M��{cO�ap�w��:��/:��* VEI��Ų�na��um����PE�E���	�J�I	�
����`(�,Q���M���-���Y��s]�����s1TI��a�be>��ЮO*Dz��y �E�[J�i;��n�*�g@BA;q?��+����ߦC��*ii�͝v|d�<�%q+�ԓ(�9`I;Ei��{��@�Y���v�	
8��޸�}�h@e�C�AA��sP?e�@;��<�SL��Kc:.�CΩ!.s����'� ������]�*~��{���s���9�T~31H���{17�N �Z�i.�x�Q
%�R~��~z�� �k��D^�0hM�7Y �F��@�N%1-{�L�y"t���	ԗ>�}ρ�%��]������Lolk]\��L����P
���33���.��mZ���C2��sy�w���>K��j>��;�|:�?e��g�J�R' 
��g��,���������V/�
e�k�Z�T��z���I�S�B�=��a��.�'�b�X��5>�84�HQ �N�R��|�gw\��eX�/��V�~��T������sqv-��J�ns�����lC�RP�TN��6:��!���4 ��EI��␹���Q�4C�_*��˟̔�I��������&�$s����O��|�N�w�������#��x��\@BG�d45�U��0NM�ݗ�\nk-�Z���:���U1sJzV~Auƨ��2�y�Pǁ��d�]��:s�����m�N�sp|& y]�K6r��򔄱�
UUr{%��=e�mErL���5�ff�Uu�P��2�42	;ʧ�
�y�k�a��xs����I�×�u��Ҿ��Oy*�B^$��ԘSȜD&>�Ρ�ro��ǁ� ��gC
���m�h�tj�wJ�W�0�ۂʁ[��b�;5;��0^R�<�� Nu9�><�R9�/�y�կX#����Q�|,DvS�:�� (Uuiy^A	}��F��@������O1�!jr�<F80K.��^�8wc0�W9t��j�ș&�8�gT�p��L���f��jd���q*�A��o���9����g�5�~���(��/��(�~���+����/��?�By���m�ܕjݑ������jq@yD���<��H�q_����1��:<���+�8��3R��s���>�U(寝V6F\I�z���P~@0��|N&��q�KX!o��i����S�:LO�Q��77MZ�}-��Y��-M��f"��    IDAT�����I��� �ih�%L{+�����
*�>� )Z��ѻޘ\��ً��U���Z�Fk}��6>%J��M�
:���{\@��C���1R��$�S*�o�2L�����
e�=�U��].�#�6���g�w %ɓxZ���Cy����O2~�����|_��:fӬ�sNa����B@��c�|'��l
|s-mA��T(>hh�QW��%��%��ζ�UUe�j�!aEe26�������oF� ���_�G���<�x�-���38 �N���=vs}�� � (���_PN{��H����J����{/���%V��E�_I�J��Q�(e���Fi�c|���R�|��d��B(*Fu���i��BHK��=�S�����I��P�0��*fw/^:P�"�:��8�☆eM�g!YI�iB�p�\S�G��@R�;=)~T)c�b5RU�F �|����H!Ĭ#ITP��i�+�C���'����@��,���[囀ƻ<�N^����K3��9��S�~f{�3�A2s:E*[ '��7j�f�q�'ڕ��)I��c;���:-����2_��_ˁL�LǢ�F�����y�"�V
�1��+ATL+���0��=�s��0j��������ދY���~� �W,|i98��^��C�l���n��\c[�;��}�b�ZV#>Z <P�? �@D�g(��;C8lD�&IZ��:Mw� ,��<�V��|Ȕb�1��y�Y�QpY�&��`�w��P9*�R(?vy��/��L>������B�����|y�h_����.�t�<�lyc8���~X��F���'ȡJ�G��b_�����c*�=��)`<?��͍^i��>�'��}���|�J����|_?'��qa�%��J��.�<i���/�O1-U��lA8'=���m�}�r)|���R٩��_��?<8ӡ�<�<�t�����pa�|{���q|Y��K�A�c��.1(�P��VJ!��a��I-+m�t���[�H+K@������nR:�s8&�U3-O8�o�$�}և��O��Z��~�'P�S��\9W,t�'"� ʏY���T'�ӟ2͙�P�7�J�u2ǘ��l}n�>׫��)I����(w��M�kɳ5���dt����8H}�B��c���̵`����*n Ɛ���o���?<�Ya�"Z�"l�G�\���r �@����CIUˡv�� �^�8*�o���)��sV*��{�&�H�E策p	K�G�R��_��ng�ַc 7�J� �<P�	��I+�9�_���#���3|�@��M��.�-����.͐�xPN�������ǁd 
���]q�!L.|�����6`�w��B�����/�o�疇��D�-l�(��_V��k}����iyP(���Oy�.���y`r�k_�?y��ܱ!����2t��H7Ojyܤ�]��iGveG�GꄤB�M�,����>s(�B)]��(ū�.��}�������k��V(r�����JŞ�$�M�$��z���O>8�G|�d9��R@�1A�@ᧃ}���%7�p&�}J�c��,�V3���K��hwg�:��ʡ
*�6I�拔ɔ$���cӧ��y6X</S�`�(/��˅<z���<@���_�����ߤE�����=fF(��T�x�2�㜃a/��b�.�=2��ťB��@��0<����4�,�����T��һ���' �h�#cOJJ��r'R6�e.c��`o�2~��	&��$�J���4�ٱ�<�Rp9�� �� ʏ*a�1���' �3���)x�>e��j��^�g/��y���^���C ��?��P^!$<�b��$��=<	P�K�3'�vO�R�9��H����G'9:(4��,��`V0�.���I�Z��\��a��c���'�`����L�ƻ<i�#���\���d��֎O��\Tx��¡|ݏ)ٶk��$m����s>�H�_�ɔh�v��Τ�"D)��L7>��#��M���b��}� �|�鏥�6}m!�|�9���
�ܡ��KI�C��w�
y����v�^�J{�lt��>�Ґ<�|K�H,�Xk�\�k4|>�p6en���{X7��\�m�N�@��H��:c4�����i(��k���(�ɀ�\:�QiE��� v�)�$ ��`�Ɯ�(E�Zş;LR�.����$M��%b�H�f�̓�`U�SV�BD��1<����2޳�J��pp�������q��c,K
�*ޓ}�B�j������b�X���^�q����s��'�	v��s�֊
�\��2��˩Gi�|;� �^yZ!�  �V�Q���V�P� ;}��(;�2;w��$���ŋ��e��R.�P(��%�"V9އ<1!�'~�_�Tl�8�:���Z���#?}��p!��%�s��	G�h���
@ʀSU`p��Յ�H��턃#�ztY|5��(��1�61�����̱�P��5D�|qƘ\���&I��P\�L��M��e����RM:��/ E@E��S��8z�2��^�G9����]	(D5�V��@��y-Y�d.c�W��o�}'�����a0(���F����@6��{5�����H����_���+��c�В J�*���bK�Ǥ2=T���f߃��ܩ�h|��P&g��zvm�*�����R��7.B��Pb0�� �+釔��+�NG�S)U��Őڟ� ���T�쀎��E�4�.��)�p�䠊�E2�	�8�\~KE���6�B�e��E��S�R�v��~O5v���yߣ26�)��L�&t�
��P�H��*P�-��ʼ��V8�#\ �u<�iF;�f�̯�s��I���Th���].�]{ 1#*?� �4Z1H���ra�j�)����5*�
���hTx��9��C���`��u�?�����\�2���I�,��ҙ��$p �C(��/+R(_S����{C��P��� 	-�20���Hʵ���d�IQ�Ф�H"�Uʲ��4'5�i(JQR]HC��&VT!^I*zc����	�b0���>V'��!fxg<��������}�׎X��ٟT��*�i��k*sQ��؁�up�Aic��j��֦�;��J��I�c��Dө6*�1��Ta�\f��T\\��2�O�ڙ��(��W�PTAA�$����s��,Aň5<7ѿ��dZ����i@+�C�G'��ªf[�ɜg�P�f�E��#Ub�2�+S@��
g��)���v:gw��!X���LU�k@�ˤ��q2".1��?��������M�� �
M���T(�v�$SC���S��ʀ�v�эh�hJF5�60f��H�T"�s�#��-��Ji8vс����	�1�J�N�"�֑��R����U{ƏrT�=N�P��}?���۶E�c������d������r�D$�O9�(N�0�/����1u��t��K��(�O�EО�V��Uc��u/\�,�*h� ��H�j�4*SK,88i����R�J�0к�j� E>g릱��޹L�&>��Zz�{�=�����\��<#)H��T���FԲ.��H[B��m�fQ�9��Ti�qa�/:�o4J���[�Rn�Ά��ǃ'|F���œ@�=
��)	Q"���,�W���Zt�� ���:����|������E�"(�l�g���k�J�h]����ɡ��ߝ#�p�h��t�?�7�|mGb�SyL�~��-M���|��Ek��TI��s�Ui�GZ�J`�ޅ�7��O\Ky|��hH�֐����"��`�U�GP����ȭh����j��i2 t���S��B��`h%��d5{�o3�7���#�kky�����|�6~=o����(���V�m@֡�cFk5��,�5�}��JC���HS���@k{r����a*���{<����Ox�������}�R��
Zk��k�m���+�V���0��5��Q�5��� ��~Ň`�Yc��  G�e�@9�"ș���y�=���ӂL�{v����^1 ��mߝ@ W&�"�`]ר��X�@������������)^�k �@��'�ɇRbBP.w��
%��G�6@�@$ a�
�1�BK`�6feK�Be�-����68�i�q{{SU������~��=޿�<��C��h���������ϟ��lpss����,��l�xxx�b��/���<no�b���o��kC�z�܎� ��C^*_����>Sc�F�h�%����4�Zx��+1Ơic����۾���P]{��8�� ���E	}U�X,h�1PZg���*�tm��w k0ǊF�$�O�t���T0Z>_U�]1r�� c��nP�5�cp �ܼ���[���ִB��ju%��Q�nnnp{{�	Ժ�aL���k��?� �tb۶���C�G�,�A2��7�>��w��1�B���x/���8		Cᄼ�<�����ߐ���:���n8�n�L�&r��Pd�&��>6ڣ�׎������B�~�'�H[SULU���
W�ר�U]����BU	���]��ANs�P�}�e?�F}?Kc���ȟd~�e�^�ɏ��0��i����em����YD0��r�������[���/P��٬����O�>��kX��e� �^ݱ��P:�?7ϔ����ʊ��j�ʙfu� )5"��RкZ�����<S��x�.�m�8ҩ1��F{: B�,pss#�KU��
D��J�U��l�a� �u܍1�>�9"���P����:Ե��|M��m]ߣ2��J)�F�[��D�Co{�}��% F`k;8���'JZ��u}3L�@jX��s'��&���*�p#�V%���^e����m%�B�O2�s'�~�Y+L�MD�b'��x�7��?����9�qL/�55����V��(˜b@�<��7��X��9P�S޹��A�r���(����b�P&+��C�+���r���fN�H"m�W���m��Y@�t�(t�www��������֮�~������
����u]c����w����P(�����������uo��}$R�~DSW��Y����>��� ��2{��c��ǯ��-uw�m�F�m����z(����>@y�'�s�	<3GJ\F��y� w?��^�G(�Y'��/+ձ�b��v�J���#F�I���|��`����b!�'.��BSͧ��kCq��AK}*K��d7��1RDZ���]*��[-�^����$ND^�(f������!x8g��d���躭��q"���^�J�8�w��G�n@Dh�͢F۵h�-�����v��;X�Bi��F�o��<��
u��܀T��!X���D���<���w��5�.����B��
�t���t���y_EO�:�ixr�˝�J)�n�?�B��#����X"WdD_�Ei��l�D������wKĿu.N���&AE�^� 0��LDP�DL�T�nA��6���Ռ���.,��,�*2�f�6)[Ŀ��8fFU�h)c��v`x4�UUGs$`�\���+,�h9�㎏�s*���aU�u� ��l��5`��{7^T��!��=�ka�9���ULpN,dM@���� �oN.�����Z�=��i\����>f!�I|�;�C2��S�~�^�f�h-9��mI������@A$�.i�Rؖ�o�OO��D䦴)5�(ͷ�E��r#�Z���B� #�um�42E2Fc�\��*t��!�N!��x/ՄR�s��:Ng�H�ZX������m�3�жb�*&"B�|I�wp��4)_�XEr�,|��[��<Z�+Wy��{�`UV)�)M� wu%EZ���6���hT;�y�m��q��<S���E��~ N3{2VK^ 囂
Q.O�#���Jk�}keO�)��	P\�$�s�M���G(��4Ե|]S/�X,�X,#x����pww�����&_���w�wx|x�u�d��Z�}��m��§�ר���z��ka]������YĭX"��F׵x||@���������{=��8�u��g$����%"�tk;{uM���{ߵI5�=o��J6��a�+�P�N4�9�MRk]kE�z��O�>��k�y�&��oPW5޽�	u]�
â�jTU���p���{l�[�:�U]a�%����:�GӂX,2Ύ�c�n�^7P�����5�s�v��m|S>5��]إ
ß�)��#���=�Y��~rP�*ݨ3*Z��o���v�La�.��?|d�U�Q��C۶PB��H�IU�^?b�]�:��Vg<�� T���m'������w���Z�MVf��H�8���{�{y���5QtUG�u�� ք��'�n7�jȕ�|�a��,v-�á�H�︚� ʳ'A��C۶�' B���n(R%$�./�>����VB+��F�X`�X�����8����-����̤�K\�8��4&-�ܺ>.�Q��&��0)���{�^���?�������t��y7~e�|�W��
{��{n|!e_�o�R�B@�u�b/-�9��[x�c����{9���B�ə8����ϻ=>NZ��PZ,#}qZ��*�VКr���Y���M��s~�C��=d�f���ݓ!`lt������"<����`�1�<=��(�b5j��VJe�����J09�<t:S��{!e_+�"7ojy�Jv䊪��b14K|P�%�Vr�پ`�*��{�z�"�e�<|pК"p��<�10Aǟ��b�Z���V��ء2Y\fgv��s�t��Q��'Z��(g*	fIY�'e�����;�1��P��P���PF�B�&@I�\!V�2tKI�� ����L	z	���(X]״�j��s=��
m�\Z��h�h��!�x��X��j�{5���A4(J+P����L������&h1R��n斩|B�C��}�5e��$�e{���2���N�@y�Iԕ)�8$N!:�������{����q"#�C1����|d7"�n0<>ޣ�@�,g-K$����|�x8Do��IZ9@�7l}�mJ��Z+x�F����K���>���-���x���9j�N�8l,Ư�r�˽1B�"Z�sa@��@yhRcǋC)v��yBh&��雘@%�m�
!	�P,�Q�FT�H� �d��"<
��`�X�)!-~�
��XJ�DA$��cf�hD���?\TS�̔�y9�P��ɖB��H��ʴBJi�%{a<+�K���I��4}�[e��v��5�&�d['�n�m۶m�l۶'פO�\��|���콮}�{=�yȐDC�q��-j��˛����@it%��YU˖(��X�(���rWsƷ����_�}w��#�M1l�X@���ӌ��4�iޒ3���)�H�T"ޖ�m9v
���h�	��k��,�҄N��F�V��*P�����H���t^I� �|�AOmǡ�)�0�[#��0�V�i�l_�a�Q�6��i��)���zRK�g�~H��Rn�D�rV '����4	��VǍ�ư�!~��p�V�H�b�l]h������N�D���r���h 8P�G�i1��~:�ö�`dP�����a���W>:�Δ�0rN�G������38Q��W�#�j�x�\x��G6�+���u!6�� v�����J$+�%^�!K�!�^,G`��Ζ��7`:���#�����Z�G��J��м#��~N�~�~��[��A�J�h����+�Ġh�8�q>x�,J:W*��G� �‟}� ���0���r�o�G3�1���L��<f��o�%p)θ���6�܌'���?�Q���{ݥ�&���O�qo�+37��\p?ђ�|���a0��Kc�*C!�z+a�(L���oω&!k��Mn�T֎�s=ܩ���0���ׯ���u�"�?@AI��S����2�&�w� �J�u���iP��#Lw�����K����E���Ͷ"�~|,���K_xݓ��=���QR��1b ��J��+�©I�����=+>���@�����F(��.@���qS'�F�S�h�)N��7w5ֶp� Ն�=��.�ͣ�w$�T'���>�&݉��0�*"���_-@�A�GIī�|��ݎ9P�9KE��N���~u'@�������DDA�c�C.T�?_��|0�{�t����1b�A�w��dz��z�ڡ
�o��eo/l8��S(%�x4U�s0��+��$\E�dE\@�u�Q 6��ᾝ���/�m���_����dsLr?fٞcq[iȴ�g2���t�,N9�I������C��[d�?_�<g$ͽJ�jk
�C�L������C��P��=����$�i��#�3W%�e�W(z>����Yf�@�ٰ��J�J f���)0�-��3����n;��5i_E���[?l	�����g��g��d-\����W�З	F{��HS9��}�C͝M���L��pm�(OcO�]*�B`�CjU�2?A�A�Nɿ*�WI�3�BK�JlDY�ms�S	�Ils#њ����H/�Mx���#C^��"A��!�K<"��2S=�+�/�R|���ʤ- 7�ә�u
��H}���$=Ϭ!��ZD %ED��rU�`x&�,���Ɯ͈�f�0��xA���c��;��.�l�O�D���{����׉]�D^I\W	C+��.w�hdK7h�m �����}��&W9W�*��h�i�܁�9u�N���t`ެ��ae\Vw�<C9�{��p	���{?&F#��mp!S�`O7�-,5��W�@T���hC����ت��pn<5�ߪJ%���/%�-Y
�����庈�ҷؾhȖ��|"$^ٴD
`)t�����a�xm
+�Q0}��2,%yR%E,<���b��WO����)�D�E�\���t����)���k�m?hT�-�4_z/ly��8�u��N������T�"&ȕ��� �L�i�<�b���m	}j;�y�=iSi2����#F�o/�O��F���f�U8@�0w(>�*Y-����������_>�0X:�ŉA���apT����h����K�,��gh>(ETz�$����/wd4�Ǻ�[.�p��h~��ʅ�����Db��s�&�[�x��� �U�ԕ�dt5s�;�S1�O2G*GGy��~�7�
-�V1pm����h��5f���_�)����$� ��rh���oB�$(idP�G�ݎ*"�}(�L-�P~ww�,%�e������/��q'5kd��F,PM���*��6LfJM�1������`�&�u��PǤZQ��7қ��e���%�kpY�G�W(������l�e�HSɫ�I�,�������&����X�N;P�F��E�OIY����f�фM�W��2�e���B@陫\����Qҁ�Lf����m�JM�)K!IaL���ٍ�B�N�w�kbʈ9��\U+�fs�҄j����ÈP�VU�ts+t�_3���t�س:��8ȟ8D��|��Z5�@T�'P& m}i�B �T���~b�z[�׼�|��eDA�q�9egi������5EA<��}}���I��D˵��̇8h�t�;_���Cx�a}�vg�K���B�5�j�eJ.�{���I����Iex��,��"��,,t]�O�:���r�N��L�Ψ����I$�9`���e�ei1���d>V,��Hj#�v�Cg����[ԑ����a��6�t.w�	c`\�kC���C�
�5{��i��3����H�p��:ׁLz���2���H��RѴ#d��S@#a;Dz�ͼ�m@l���h��u Ʈ����o��a����{�z'�	]��J4�PD{2���s0���P�$c�mK-��-mk6��24�Y'����}��f����sy�S���1���dA-������� ncP�Z�Q3�&DH��1%��ژTiS�O��\1�%"KH���*��Y�_jb���Gf{8]��5�U��.~�{=(|��|�F֢�	��˒xJݶ��ƓD������(n�SY�*f�v�A�W�N����2E�K�֥�d��&2�[YaP%!1h�����~��{~����c�aE�	�U����"��l�|a�3N%|�$$؁��A�������av҄:>�ܗ�Wѹ�1V�ڏ����,bR�����@\�5�I�1r�<�c�+o�=/(c�NHb�F$�ɥ[8=���1�`9��;:�xH�k�M���n���\�~����$[�AC��	RZ��Y�-Q�ɻ��RU�����=u;Ap�Bjj�]}c�C��O���>>��]WYq��
\q�.�h�E�~�Jӓ{u%�I�9D#����77񍨏��`�n�e+r�w�,��7_�.^l�c1�@�;��lN��84���$�}��=yK�c��9���M��Vr���vl���;$d<&ϰJh0����(R[^�F�쳾X折f�F�b�L�5)L�M����ZEE��N4�m�P�Ъ�w��~�X�����Lf�����6�QΠ^�U*i`�w&�]�u�;�sd�G=�ø����k9�����%Frj�1��o�mE#���X��!0����Y��L��S�� H����̏���&��k�3�X�i�#����BQ���Cm4��-i03�ĦA<���	 ��M� ��(�9p�X���q��dV�0s�n��Z��ˀ����t�:th��-���c�rM���ٵ��f��.�Y�*;\�^���#q�H�2��%L`p�{��g�V6<�G5Q�������sf���!���+�5����\{�_p|���Ry�����k������q��[�\��aץ��Z��#�����H%��;�I,����/
g+��t�2-
�t���ZiLz�9���ã�ک����DHL�|��U�D��z)�f��Bu�T�(�+Lٜ�U;�?Φm7�+ߨ?�� ��a�`��i����Ԉe�;������\/��fܶ��!��\�@�U5�����QÎ���s�@H�LO˼��Y J�lU�XӰ�'E��2|�2�����bg���(0�{�jX/�G��m~�`�z�����}[�ٷ(�����ʢ\�,��H<�����%e��I5J��
��j�$�&�u�C:�E �Xu�eᏽ���"�)bA�c������'}��o�]�{$)��T*�ADD���E�q���(�m!kQlQ�.qXH]��;|s
�����*�Q�\āL�3|���Y�1�2愈�S?+N�\�+���\���R;Y����� epe%Ձb�V]��V�A���l�Ա����_�`ߔ?z"E0_v���_w�'�����`�Ǖ�a88�&�Ñ~Ceu��p��b��'ѝp�^�׮;~<���}���IU���£$�xPtbëI�}�Cz�&9a҅0$≅#����C�f�;���E"v��+��r���]SU`�^�O¹>��u&����0;[E���{;�u���>���q�VM�	}BǱ�.	����e��J�;�$HBU�����|V�~��5�qJ�o�p�B�2���0��X�"a[v<E:d,y��m�T?Tr�{f*�{O�4�)gjH�\�}�ǣ�肏ڐ�xG|E�{z��^H���Jc��]�8$a��?9��Ƞ`O����vE�1m������GmGj�+(D�,�7Є��˹��ۅܢ�NfM� ���_�EFA��{'|޿���%		 �H����/����W�d��dH�n��.Ɣ55ZA��V�wR;�kS�A���;�*<+�W�!�UR�1�@����3�n�f�������N�7a�����z���HT�Z�E�q0J�ɟ[c��w�=���!���:���yF��$!�L��9��(	����թ�p�`�']�7�������"�܉n��>�H�Ҫ(�A�x)]]�6m?�`�}��M���U )^nɠCǨ#嶥�\�0+��7@U�Z"����3��#��E�s60�B/����:L�牷�������	��^�1�3Ï4�n��rCP�wt���O@l�3�nm�-������Tyq��KwKze�ʬ�y�!A٢�o��*SYX��NT�Bk��fcj��������-ٹv1�������� F��vٕl5�do�v+h|��w���'�+s�:�\*��ʈ�����-�W�(�C�O��s\�و�[x��Ac����^P�M���O+�_ 9$�ꘄ�A+*�����#�#
If��Eyx3m[kpd�����!}�Ķl�=»�JX�k��.�P�xjjCڼ�SR�&��(h� i��k��8}�7|�/f�Ċ=z���[*@�r����K���%x��r�B��h�h�/�fn:��՟C� ����H�
 #��3�x��2��DV-��gC���Qɴ �'���VһFd�b����fgb#�uD�K��7$�y�H��N8 �$��Πg<xT��`>7��h%Q^]�MCno
���|Q�)x7���pf]o�n*hB��l� ܂��!NL?5�l�c"ӠՠKឞ��[CQ�e��S���]�+��fE�|:	��<c��/�>)޸mz\$|���M�I{������� 4�DZ�{�O��K�w�/躝�)t�% ��<�͚f���!I)C:��R�dx�,�m���PR�� ��K�@���X�&�ko0B_�Ӫ��� 烟��@R�-؀7p�mek��k��'���B�0�[�|�nC�ns�srOn�Ȓ��~2?������۶g�VΩD���Er�x��k�8~�bڑ�v6�&Lr�Ksk`�!?�(���(����w�{w��f4��0�R� ���C�&��洺{�f�@��j�B�Y�"�!��z�?j��Ъ=����_S�76_�pT��u��£�@F$�4ا��'�G�=+ӥ��u�-l�}���Ut`�����8��Q�s̈�-� g��/3�5�T�B	��np����t��Ay���^�pN ���i�(�?ȫZl0�RS�->7��C��O�ѝ� ���N�p5�>.J+z�������]4�,�e5�[���"[\��J����$[�ۦ�D~�y#q�MrY���z�Z�Z�Oִ�OσZ3R��U��ã8�o�78��o�(|��LI����<��*gL���w���{>C�hԡXx�m<�&��
�d'�G�E����[mس��kqU�iXw�]�Ŗ�O��j���E�졙y�A1t�H�þ����}ā�� ���_��im�z	#E��/�+[�
o�b��0� ��a�?�K'6���N`�Qk�9��\�4��SIJ��ǚ�}��5WQ��q'�s���*�I�sd��,k�%�W��ĵ�ܑsL��tD,�LJ�I��h��c+�TO}����I��Zj\�"%3�U\��*��E�Y@GB(&�gFcr�S*�K�ʉ%U
�^��G��j+�}�LB��"��;4��ϧ�Ž$��>��rW��\g�{���.v��й"�����qrܣ���к�BJ���9D6i艁�q� ��S(	�w�\�%UG�G�Hd9ˀa1���yi,���"��#v�-x틅'�3��i�x�5/8R"#�GT�n}�iY!du�[,ѱ�4P�~�a���=��$
@e0�����:���^U�!��͕M�L0�CѤ���G@��F��1�5�2 gI��
�� 	ۤɉ^�/��Ҝ�5��\íj�
�;��qV�D$�6W��[��<x��8v�$��y#�>kx�����Kj6�x��΄Lq\�ٸUy|+ �a윮�,o������|��Ǎ�^�C��t��+��n�IV�m�g#�#�}��k
%e~��+��':2%¬��Y@h�T�E�1��
�赇�q���@Ǉ9!謅F+����զ�G����l�53�f4㮨��o~��}���7�8{��r�u�%j��<��)cQ���Y�{�;��%4
K��1�+�[����Uձ�Sp�%
 � ���b�N��Ϋ���%^�#x�$�]�V�u�Ü��`�3O��Ȩ��J�L�ͪ�)����*4��:Eo�����,����<0u���Nj�0+�����t�[Î%]L�g���E�����V�	�f�^��"���"�!�q�I�r��YZtHK	�
���U�+�L�{�n����+��?Ŵ)�������! X.�O�'G1'���V�-C��
k�]���&��&M3�4��E�SCV���|�}�W41xY���� u��������$�oD�`�i��R��~���(���t���8U��2�����QpxSL���cY�������ߗ	p�N�U +�82ӓ��Й/)��rx|U:�f�ud��̞|:���2��yDX��@,H�����	�����b�D���|�-򿶛= �0�Jm�I>$��Hm6Wv�Oc�zE�wk�fp�O���ґj��V���������޴eR(�� ���S�6���Ё�t��6��ڮ=lY���Q����丂��.�=��VVgv�^ȧA;��B(`b�3X�#��P#��eL�2�	[� �a�[�4���-��L�e"��@f,���=K�y��^�#�eAG`p�o����\^"��KG��:��x½|{�bܺF��ޙ��0��A^]�Y��[XUת;��?	�m��5��[�&$0c��o$��-�2B��
o��'-,��i���'�cS���ܠ]��C-2�+�jX^�^��qO]C���C��08�������V��I��8�"s4AH��"K���h�ޱ!������'�@��H�<�kB��ڪ���_/voǈ����?h�ޥ�,�+<_��*�����֝�"o�`���o���}��=���Ŷ��W"�e��ӟ�i���G�������3����ȬiԬ)̝�5��k��S��YPa���AN������L/��W{B�q�j6KMŬ������);}0�0Z4W��_�	$����`�SAxU��)�����r=QK�H�1
���u� :�*M,����N�p�(%d�=u��z�sI�F//�utuMq�Va4�h��z؍PGb���uj����+��H�w��~��������c,U�pX��69��l�*q;6��tY��妎��0��0�Oګ�&�s�wY��/�@�~���\`-�� ���	��;u7���1������3�F�%���}r���&k}:�X����5M�{��+e1Ls&֫�k%5̝>��=�bWn���s<���x"��������e�]�h3���C�~�bZ:,�?=%(a:n�F:��}� u/֯ �ZD��4�!k��*.5�]j*c?r&!d�$6�$������������a����U�L@.��N����7/}��[#��7g�DK\�F_z<a�ԩ����o�HQ x&�7�c �#�����NRm���i(��R\�����O�V��N����{�I�+*!˲��БJY|IW��B`5A��I�y��VC3�VӶ�p'7 ���`xK�(?�A+uu/�]��2l=̻1��������?%�:5cHhS�U�G�[l����	.��F`��fg�(�[<z��]�sI(¸�7]}-�΢f���/8���%������Ƨݿ��#C6a�8�A��?�'������r�'�����e���a/N5|Q�y_�%m���$��ܽ�W<�HN��e�&�Dݴ�xL�}_j�I�Y���! ���<���y�_�)��6jF;� ���iyMq��MԑO������N��Ã�oWlq㮞1��'�-�]�;���~�g�!����,X������)�|'����w��J���y�^<�����Φ��il�8�Σ;V&�g�Z��E$����[5W;H��Yad�t:�QbQ��y�f4�՗�[�EU*	̳�G�/`�w���^�o�:��+���6h��X�R���~Y�Y�Wm*�5���G_Y�n������!����An��_�#����j��A!�}ZKw�O$�[�1�}������w�v7�+���I!շ���/�DC�L��w���V=��I�׾�z�
f�Y�j�bw�ۘ��ơf$9k*āŗ���t�t6#}4�bD*�B�@k���~�����E]��߿��=c3�=�̤��W`۰!`Ԡ�'�]Vi�jI��:����v�cd_�ѰQ���3 `lL��U���c��Ob��@�j)�J]������H�+A0��L"ѯ2+K  ����]&"�DF����He��a�!2���>����͵Kj��MD�B��;�F�Ź����QmK1�$M^�.�F����v�$5��ʒ���;��A�@�B�ͳG�����%��.�Te��fo��	n!Dw�v����|��Dq�O��a��Y��h��W��������z!�Ƿ��E�-��`���n K�����螃���(d7 �Ȟ8�یD����tB�$G̕�J�Q^��ݨ��[�]�v���'oʗ��;����}
��^f�F:���������,��Y���6[GZu�v?�R���ZM=�B_>��V����_A%��}����Mi�����;��������w��v?����{��urr/|�����ׯ,�^"5�U�x��X׉è牡1�}�z�PН���H��y鐿1?�};zVt�~݆s݆c#c3y�I�p�C�r�S�6� �W�F��;�2B��V@�vT&*��4N0��IІ�/akR���%WD�������_��ޡ1��v�(D��`\k� D�40��Np40�P�#��WP��Fّ���%����`����������8hG�9D�
ƙE��b��$��J+G��/#.���#v��oZ.��.�E멷����Ynx���g.a,��~�ɋvD���R��[2R]����o9���uR��0�j�o`Ŝ�������_�zx{Sд'�m��������Z��U ؅�u��խ��ܟ;�����k��?������v`]׽9�`�Wb����	�@�����vP�(�� +c�aZ�	��E�)��eI�岪ӓ}g:��#jȌ�`�g���p��c��;8��KxD`��O�m�i,���-���q�ۮw��8-� ��^o���0��gA��g���Qo�R��cHi��Te@
~�:q�K�32<�x�����VE`�r(ר�m����)�7���|C��^#���n�����s/ؤF�xȍ�m��\Uu?,B�*����\hY%jИ�Gy���!�0'yԺF��X�ƥ�������0�oCv\�a����#�=���F"���s;�6ItZF�+ӿ~ d��Dm���=��`b ��dh�GI@P��ޥ����8˺$Ԏ������>�'�ύ4��TD�Q�+���O�:�la�
��n���y�?|��ʽ��cM���:��52~$D
3�4*�@8\AY���Z��]���C��]TsB89����/��
6p��=��EV�5(��5r �����3��O�5�S3Iw�tX��Z_B)�gf��?����q�(xu��%��-�N���*�,�9�9�i��.d1�2�ي#c�{���GP,���vd����W ���{D�Xa�,�ҥ#�:��H́I�1�WG��<Y蛣��@��ΖRŲnd�!�����o�6Fډ)<ͪ|s෱�1�8�٫�L�ߑ�6�dҜ�"{�")�� ��R%�?�o0�6,F�]Zß�g�r]�v�v�1��B;��[&ɮ����y���b`E����CS��L����k��XZ9��}^������kضkذ�߰���������%�?��O<����b���s>�I�<��`Oy�Т�5�P&�t4"�``,�	�@'&������
|t� U)�ܢ��:c��ȢZB��#6��pV��sZ��W{�����z�U׷���bӶ~����̂uŨ��~&��_�l:#��pV>S����q�>��]43z$MS"�v1��=z�7>�ֹ"yU���Q6륻����HCJz�	y15��c'j�����P�Vk	�e�b�������l�B���y�h��?/��]VTj��^{���2��z��G�J�]�b�1��U��O4�0N�,d�:@�Z�>A�Ժ���dVb��t*��G� 	,�J��s�R�U�3�Bf�R�rؾ��c�����@f��ڱ�
a8ͺ5��/{Sh�����(y:��$�k�>e�;�9|Ǝ��N�A@�ke��IAH��8㍿�����M��k�vk �gip�A��l�E ����Ά0��ߵ��K�G��V��t��3�ꍣR\�_�f���k��R���
�1���|������H������RG!�iВ�u�;���6�V�xp֚\����%�9zb(O��R�7Pfq-Ρ�|n�(	a�V!��o�]�0��O<y�0|I(���1 ε� רʿ�B�G�]�Ě��Q^��o����;$����%���7ur��'��:�q���.a�mL
�2��(����S[��ûZ��p�8u�Am.�md�Y���v�>�)������=f����7-��X!�o��k�D��_�}�v��a�=�(}�IK[�L��7J	�o�B��.�>;��<�7���4G3R
���i��`g��|Yx�C�bMx%���y\S��s�����_��&''' ����1������ �T���C��(�8��k^�y�y�A1��	-�̷�N�>&S���pd?h�!˘��%�a4!�E��XRT�-�����]�t�#!^�<�=>s��j3����]���;s��[�4[,n����{.����o�-<���+/��#r�#���=�N�#{۝�.�y&�6
*�]y��7��D�1*L���q�W0���B�/" �m�a5�+*^9abҎM�t�h��	���2ʏnȟ�9� �ų;�b��AcE�=��;.Tww��0����p>�}�:��*������qD�Y"��ڹ�,'�l�\��A�/o��&]z�Φl�t|���O�ķX�ڲH�Jxⶈ�Vh��ZX�^�_���~W��W����x�j�t�qN��P���^*�^m׆��Ȯ"�7��MD��(Y�(ᎆ\�J���g����lu�P�"���3����)�����L!��͠�fq��������=E�0L�ҧLsjn��}���v�'�>�b�p\����Ї3\��d@4Pi��+�aV��#�/��㟝��Np$����_Z�lY��u"�`�7';9���)Q�X���/6݇c7g|oɐ����Y�V���	MnL&�ܓ��<�_��O7p
$BU��98l��[њm�,�}j��`=|�7׬QgRsu>)Q�<����Ct
C��yRZs?�-���O�`�J�.�Q�]������U���ͦ��Ԡ���}
Fʯ���/1l)�+���檙�cС-D���]v^d^d�Y"�ĕp6��V()1�A���W[W����b�� �����-���TKv�h>���8	Y����cM��� �ę�̪9��ٞ�J��U5L�r{��c{�����ϩ�xo/E�#�3_�E�☫�Z�[݀�d{�2�2g�g($C��l��	��݀���
j�q4	j�8�=����l�4�6�9�p{�3I?�wYN��6�*c�ЩJ됅0]���`=���<��d1)�P� Bb9s$w��6����3��C9iγ]�;����_p����S�W��)C�1
w,[k�tU-�A �֍���E�'}�<>(�I�[0�/�<3�f���S ����j훴������~R���@eԭU����@�������ٵ-���,7��M�^��-y�$����o$��'���(��;�2�3�7�d��M��~���D������Ф��;99�oo�I�V���j�����T�*
�.�����E��7Ј~V�^�!� ����@ã�Vx�C�$e�vC	R�Z"izx00��9ǌ�>�9��#:���N�RN�QM�(��!���h�N^�֌�����?��}����3��U�S�����G��ۇ����<_��.q=`>tO,�J��mk� ���阮L��%*�3��q)B�A�4�3I�0>Qks�n�n��8E�^MLE�j��O�:::Gs�Ye�"�1���^�LK� g'�B�� ��z
x�XHT��  n)W;���T$+��Wan���(.B$ȕJ�&-阇K�e�7۞Mz�R�a��8��:��M|
�
R�^1���?����,��Ӟ������ܵ�u�}]�{-܊P�aF�Gl�Л��"���3�5bу:�&�T��W��%db��չ�MVɵ��.	"�tg���0GVI�~ЕPX�/���j1Aݛh�i�;�Z�^��X#!v@�p�.T��{�ϗ��+�jE�����}��A�ݺ�e9�{{	q[�4׾]��D����;��Bv��:�d	�6�`���gj�w�F��Z��C��qS!����3ޕS*���R
`[F�����ˊY�O��վY�Q�d1�H�?��Q�L���|w���ܬ_���_������j�n�2a�}����9��!��`�����u��=�G�w����;��7[����Hh\�67d+E�-���hH���<�PzX��,JdW�ފ�֨�Ob�9����+}�;�.aqҾ�IQȍ��ll��]0���v(<��:�&���'B���Q�q.Ql�\naj���./��Z�r�$�(���f)ҵ_k8|�XӤW@�0��=���G �}�Q_(������:'������P�Uo2��.x�.zۏ,��q $��Î����6�˽�ʳi&�%��/��!x�׌�)�v,�.R�l��w1�t��ٞ�,g
��lX�ߜ�b;D�l�,3H���&�QUtIɁ��N�r��n z��K�_x���	�n�xץ�Zڜ����%sM��uu��Y��n�ٻ�s���݃���u�����Vo�5�D_��;~�	��__9�ֈ|I���4}����<���(o�YRIX��M<+���Q�� �&��U�?s`��P:M�F�21[|��uR��=��W^���$aW]t�TO0 ҥ�p���Et�i�$upr2;��*�Mm�f�����6�&CzE6�Z3�4x��U͐�)T��x���Z7t���vo��N��_F�ϵm�dK�t��dg��9q�2�M�����N�s˖ R��	ߠ����Y-rLU����x4$��%�/����������-L�)»?=!Ļ�;b���;N�8H`"�)Me������c*o^W���i� wX��}���pŚ���Kȹ�jdEa�T[��MJ�kXy���x��
LE�Lf�lec'X"�,1����o����+C�FӁ�cb	nʔά$4cs�x���G�i"m%;�8#X w����
����Z
��>�uRK���-*$�1GaI��a�f�e���Ӣq�58)[KB~N��W��Q���>�PF;�WȋN��b�5�ju�8�1�Ԫ����������D��*Ѫ�
�CN��@30�9zz"_����;c��b�`��������x#��,.��L���z�U"�CZ���{"���o��>�:�M�V��׍H����3������,�6�F�p�Ҝa�{N����xU+R�5��]nP8��{_8�8���Jg
�P���b0���fx�H��	�_rp	
��@��2|7j$B����D�"O���t���G��sJO8N�$��oB{�܌�8���q�I���=@�x�	�ߵO�
�阈 'Oԓ4���s'��~='Q)�-H�rEv�J�=d��ѐ�{6���<�nqA���l��R�%3��%B2��hmy���/�n����sr�-l�|�Sl�3*�j����igO����~����_�خ���a��O��bIՀU����'��NFsݻK�߭w�`� G�Z�ɪ�bF��A"��nɺ�$a:#Kj�o�fl �0_y�j�Ƞg���Ġ���1�̖[�	_�9���[ T�Iw 
�j�4�%���M�ZEʀUK��W���[G���^���5��	aW���U���L,9	�,\��A���:�#H5���OwN�񥜁�N�[#�
�!�af��X�� ���V��+�۹�"RtZ�xe�	��^G�qA܁����fG�m�5��^Kl�ti7&[_�QSAN*�*����쨽 lBeb��W?$~�^�j/ o]2Xg5�a�����x#\m]�jEWm�Fl��J<P����ܻv��>�O��F|Ȱ�B����<qs�K���d���yR�5vb����/�(!��%��9iIB��Z|60�n�rDV��-��3��)��[�/C�t⊕��W԰{���%��� �L=Bښ�m��ӆ�K�����F�Y����E�IJ���a�>L��!OZ^(��S&H&�,<W�B��Ǿ�놭ˢ�����[:�I�;��Y����۶���E��cGI����C�1ea�!Յ�� �L�5Wn)�
�����X�Y �
nסSd��g������J��w��^��q�;y�̺FVV0ݺ�_{S�r�`Hw��A��`2˯�˄,sK-�o�Q+V܍a����J�����T� �ft�$[J{�����B�!�)�,#� ~�J��B>�4����<4�տ��a��+�Z�x�N Rl�"��ӂ�J��3��cD�(���m�m�k��e55�,ӣx�e�ﮪV:���[-Y^�ꧫ�9�흝Q�����6X�h��������ۿ��~�q���~�����3I�B�.n�bKl�d���('G���oȳZ��tO����@��e�#ݼ�IeʝQw	��Sm��U�S\����Ռ.���i�ؗq���&���&�x���st8�9 ���	 ���~�P@S)��>QvZ"�աvȯ�1,j�5�4�a5�&��e�ҫ� ���2��7�s��^Α�ќ��?fw�g�n�SS:��n?�v�侳&�9U�@�]{O�g�{��g�k��J@)��Np�
dE~��԰	�d�n��T���*�f��c�����)�$'�{�E�4O����%��������3��[����z6��l��!@z�O���5�@g�~$]^�Kt��XHu��e��"�rfjT6���~Z�;�����y���^HB�G{��a8��q⃨����ܐ��@X��Q���V�YX�u���;��������ﶩ"�{@B���cH"ysO8j��I����g��'g[K�V ���o�pH*R�t~��L�GYǠ��LZW㱂�T�תuȈ7�����K�a%��e^�l]�~Z|Y���t��p�.��{�����U���� ��4���AK�Ԥ�E=�@�1�?Q /!Y�$GD̍a��R�m�R�!O��<&���12���=��{�i W��.wy��}�Ɨ�Rʺ�M�?RJ2�� ���B\�&o<( �#V�ȃ ��l 80T�S��V4!�����9b�¯�9!t�aA��{��f���c�f����4%V{xE�C�Dp�r��?��i�� �@:�[R�Q�5�M3���x�P>yP��o" �&W������-$�=�W�X�/ibe�5#Z�8Q�Y�#)�s7Pe^�M!11D9�r	r���X�hA�b�Z+#>C�$p��OG��" J�3wgc�<� GM�|�3XI�<IZ�a<���0U5
*t����!l��1C�T �Qpn�¦����y���
��)�
s�$N���99/4��TfQJ&D�!?�����Tj��S�\ϛH�+���{��l�P��S�u<��3��s�Sv;hrR�E#eLUJ(���>|_C���,a��P�MJ����Z�+���8)|7E�x���_U��tyƲ�DZt0�"-G%�G�El�Z+�U���D��n~��Cbz��i���P��`���'fVE��#�_W2��b���=zk�l�u���Ԩ�LQ�>��.k�$v)��<p�sh�����(���n@��������K��1s6������6����ģj���(C�z݉�ɆtOO^�L���X��H�F�5(�,�Q�lu1tB!Ɂ-    IDATK80�%T�x��a8 ��d�s~�P\b�*��py/P ������A��{�9�'0H����jhS 8/��{.�u�V)�y�{��sr8cG7IB�5�p	�{\��V)kM88NRՓ�P]L�"ú��5��͟'������x,y>50;����$%:��������X���}��<�S�Q�"�T�Yt3.c�{Oq�B�0=���J�9�ƶ07	�0�Υ��������P�`�0�u���[�CvR\sY
�R���P�brY2d-����������B����_����'�������SG��f�˖ȒM^��ϒ�`�'	q�c��b}��?�@��8��l�A�yA'����N�F�&@S��\�d���Vug-���+fr���I�Dt�9�J���� P��M�);K�iWI�����~O������#�x/'��~^�x����c@y�"\,,�����OmWC

UV.w΁�fk~��5�� # H���)y�`ڤ�1d����� �])�
Z���H�_�48�PE��d���嗚e*�dz?���vҚ�*�Yk���TiXke"���d	�^>�<�&�D�� ���A��'
�H�Fi� J0�b�sL&'Gl��Z����(05���� ����dg�������	Z+(���ܮ���-|@�����X�B�Lh��e?��AS`��GJf�<$WX�NJ�Q9k-��PZ�C��E=�HVU�z��|��Ozv�t�,�4��m�4��&/����.���5�,�wq����`k�҅N-O΃m4�hKT@#E���� ł�4M��j���gON�Z-Ez�Z������#>40�%�͕><��G����1�&�ő���y����P*�F��9A��9�|�$�:�`�^����;�:�P`�r��c\��s���HN<�Du-�;��
��)�EiW�rf����I������4*%�J9��� ��*v�sT�gF]5��Ev4T$��M�³�/��������ϟ�9�6R�{�V�ZLA��2���t/�o��떌�.�h�f�F沞��J��4���a�K�Q��ʭQ�d�2��uc�z_���H�H�� �!�W*Sc�, "�J~�v=��a)x(�E�j�0ٌ|������a3��L3��DrP4l�p)�	��gggx��9^�~��߽�w߽�>�m���~�O�KD\� ^�@��k��I�x�nl�cz(�0(���n|��	� Q��$+��*���)��<��;�2x����|nl%$�h��e��ё1�dI)�p΋і�y� ��77��8���
͏@���4s�	.&ys0�n��Hɣu����&��=y����������Wx��)��,x�PU5�>{���^�y�bp���}�mtχ�1�ɍ����"LL��p�(B��0��015�SE�[�X��c�����=�ϊ�����O)�q(��Q�QJ	�5�ޡ����Y��?K�|4�H(�ͽ,�B�c�X3�uj��BeTf��Y����F���=���?�嫗8=]�i8�q[0˜�uɖy@rf�	���y�@~ ah��<��XWv�]=��#���ܔ�$��.A�q0����G�p�Lhb�;`���1�|�Rh�6ƀ�x	��YP83��E]�X,�rbq@�7�m��n���FS�9��B0�����|YS�4
Z�:��]�V�F]/�h�x��%�>{�ŢA�X�ի�����X�����j���m���s��?���~���&{9ߌ�L�����0��0l�� 6tu�A@I n��t2i2*�����}E�����g�����&�_�0���)�����3ɩ�{l�[T��sVX���;'�r�D����I�s�2RRDg�b_�b��h�(� %8OU-Q�+,�S�������x��;,�,K<{�/_�@WW�h�����6����v�=���r%2�4L��|��S�����4�5)0��$�o���s2�3r��%�R�r$�\eK�;��w(u�[~$�=8V��ttd��L��r4���la�����*�%�U��	�����y�)	��T� �`�P�a�9��4"��t�iX`���1�^�jy��/_��ӗX.N�\�q�>���t�0�y��� �'O����3�}����d}���x�`m7���m^����4b��Y�Ax���V�������=�Mbj8[6�!HM�7� T���� PU&:06�����lV\!=���L��k�,}T�g�[�)��̰������c@y��R�B$�m�;b�G?�C�B@�w�n��/�$+�*o��r����e)��^*[�A!P q�V�q����D���u�YU���'���
D�'O����	���h�U�N*(�ὈR� i���pgg���*�8N4e�K��vDS�[��P��O.>��U4fO��(*D2��d!
DMq�� 5'�D��39�R�-��ɿ3���)Y�`dZ�'�@��"�rJ@�荭��U����thE2�����4�r��3�ω�(C�$����Ds�b��0x�0�m�/�Z�pv�}ߡ�;����u�<K��Ik�
��pփ`�`�JqN$����j�'gu�4��u����~�~�{|���ж}�&��.�u�s��m�u-���v����%���a�ݠ��a������[�i�.���\('�m��B:�f[��5�Bhi��K.�H���] 9���c@�\E|��[`r��D�����S�$�h����=�3b�uyy�'�C� �6�1�����N�(�P�!Ʉʞ,O���s(%�Ƌ�'�5~��?����x��w��7x��]~/)�^X����������v����
��n7��n���Y��Bi�.�2c%�^�����Q�uk샊�U���1�<�G}��)������{��1�Gou�r��9�������@E-Y"m�%�}ۂC��~�8Wb��z8�c�^��FU5h�^�x�ׯ���U�V$������ 3�͛wxw~!iy�2$h��`{�P�v�n���6�tP�����Y�����k��
yl`����w�?��ʑ�9R���tr�[�*�I3or�($7�ݝ4ӓp������s83�S�jnV��s{��������_�������3��#���.�EE�a���:�ؤ(�~�r�{E>�*VU�&����:�����<_�h�Z��}T�/Aз��X�O���+��w�15
}�c�oB�����=޽{�˫��������h����v���c��E�6�+l�װ}����o`���Ǿ��졢2��#�@���F�1����/R�����n���]iK�l#?t����/^��C�TAe�
S���X<O$���N�2����J�$�rhO!�Hh��QE����pr��:Y��},�:��=�v�ݩd7��2���j"��{�U����4K��>A۶b��c���rѠ�E$�H4��Ԣ���w�6�kl���n������H09r��G	�0}G���O��;�)��ݟ<lGw��������d�Mɺ8E9;�1T�Cq���3�g8 e0[�!x�O��W2��R��MgdC%�#�>�˽��)-r FC��Tq�I&<�,�X�6��ju�Ţ���Ǿ�c����۷��C�@�.OA/NVx��5����������'��ß��O?⧟~�j����������^<z�1�wRc��T�5�&�m���UB�~���K\__��Rp�Q��W�Y��ޣq�7j�����㚳�qPI�=w��)3�,��?��!@���������nl���E ������D�+h���A�C�B��m>M�*��xo�,��D��b��bk=����'E{��b������4��r��>��K�f���9��ʀT�)���6�v��p���
�簽�ھ�v{�}���{xg�.K�ؒ�!�ga�1�1j������g��G� ǂb9(�q�0�9��N
*�l��*���s���]�q���{`M��1�<t�yp�Ҡ�*�
JE+&��ߠd	*��+�oat����u��6h�
�E9�FK�$��M�$�\��b�YUX.V�ʈ��R��}������������oA�4 EX,T���~�M�շ�-���V0��z{���s��DUvi��(��d�g_�<�g>�&,���H�t8p
t�(P3��:<���&����SU�x=@��?G��c@yP�DF���.O,�'�q�? ��03���EEe,�kP�4���1���-$���	NO-���]Hi#��M�䙡��ж-��-��X�O 0../"��Z����xw�?��#��EߵQ��`�����D�_.�P��v	!�G�@M<�oB�d'���8V��|e������7d �*|)�q��GF��ޣ�L"���pk ��g��z7St3��+0�ʧeǵ� ]�CT}PZ�2d�&�n��e��4(��X,�X,�5�i�D������ZΫ�'�a������(���= `�h���~��f���W/���K\]]�������ڀ�~�˫l�Whۭ����&!��d��aL�Rb�ŵ�uE{�J�O�V��&S@r��Y�����G�8�]��`�+� �F"�y�b���M�d�Diu�:���m��G��1��N�!3��J�>�߰��h
�"����A�_oE�U���S)d��L��ފ�=M#M]7x��)^�xf���5����C!�O6M��ϟ����y���~�8���
���l����ܥb�절�	P�#��jp2L݊җ�P��'{R�&G����i��t*�=K��h������R��IN��� ��C���������O=xR��He
~�:?��2Y��Ǳx�y<vy>mogr�L�3�I]Q�����|.�	F����f{�E�x}r��b%��nb����.�C'�B�����d_ ��v���r����	Bp������\�mwh�o��k��ڽ������E�@yk�ڣ�V+!e�AJ%��G:;w�S&N`ԙ�.�x��.e�m�b.�����c�NΠ';X�&������Z�"�"(�w�Ǉ `I��1�|��"�d9[�Pd1a���l2f�E�ڶ�|����0��uS�1��^60œE��X.89YI��w��x��k�|�?�����_�M�\]]���7��w�$�^\��������ɬ�s�\�R�!qp�'&bs]����.gh��P�i���������{����ʁV�>p�L�2�>��e��!���1����J�<�I�DwGcd�5�G���L�~��� i3�GP����c�=Q�U�<�\�Ȃb���H�`��B�yA��-.//��~�Ø�xS��*�N�rIE�$#��mquu��o��y���]L�k8o�!�G�2�E櫍AU�Y�#u-��g����妒��kah����Ld6)mp4{aFvL�NO� �K�,�#���o	���%
�(y�C�
f�F�\�8�Ǆ%	LZi�жB�o�M����Z�X�NP����t�qQH��� �ʀY���
o޼�!
 ��AD��w���ߕ7��MEȵ�N<�i�p0� �I7|�������ñ����-�q'�
)%-�>P�5-�\��mcV��=0n�Cq	��,h��{(�E7C�~�|�U��ѓ���y�M����P�W �D	U��t}��n�,�g*����"��5HI�J��R
hf�'�����Gl�l78oa��D�^�
�2��1P*SAi�D1"�I���������"Ok�-���O?ٴ`��'���IY�$��FV��>�8����lf��3���3���j�5*�b�U]�!@��Ѷm���,�%O,'�m ��8���
	�3���zu��ۏ��g(�3�=;����0ZHH�5�Y\��e�fY\:c>0�e� &E1$E�f��O���k���������S���u�����#@�h�aJ�Yl��a�\����_�O�G\o6�:K��U�h�Ǯ�@d`���Jю�2�7�E���<�l�Ҵk����&�y�� &��q�vd�~�~?pX�_�;G�l��0�*'���V4t|�BS7 �֏��epS�RK9)�m���EqqE�USp��i С���jh��}%��+����( C�����/��E���eT�i1
���gY�V�TU�D�KT�,u������Y�p�N=����\
=�;��u��0<�J/��%&�8*��L%�8qo�	�E*���V�%%/\���@t��i��狘Y
(�<���њ�B��9�z9��|ރ$g���G|��K#�s�f1)fZ�8[G��x,y>S������BSԇ�l�ѯ�,)�Ve�𗜔u�D^I����i0F��A+C�C���9�M��n����y��@�5�sZi��� �s�m��oἅ6��n��농 �wH7mt�guY����s?A�Azw#��8ňp���<F7C~S�A&�����^494$Ԕ}��U*�ϟ�J�ʂ@�X��y�M�R>�!Z,�<ȗ����u-��F%BG]+)��`a;fN��ً'�B�T�{TUNOO�X,"��aߊ�c�w�V,AZ:���0w�RP��.�-T�(geC�����������]���u>�X�<~�q��Ci��A(��ASvN��T��23&b�
���� ���|�\�X94��<��gN(�Hj0��a�L/��\Kw]�6�-���45����=��f"�tz�\gWU��h��6��BQ��Y�Ŕ�D7�k�;���Z���^29��hy ����.n�/�-g�: q��I�F���~���1����&q�����Ǌ�+u�@�����P)|H���mLwY���JYM��TJǀRc�\��d%]ّ���~���VD�|ۧ��am���h�1&�����G�k]7X4TU�y*]�b�Y"M]��KL�hm�{InvZ�h%���(>���q�rO,Y:�R�<��
�MGG�n���yA����#��A�7��"[��@*�O�GM����YJ�'�E��Z ��b���sK��+,�K��l�x2T����}c�[�z����t�@Z�_�>�"=��5@[��gRU{04H��z�����a�\b�!��w�8??�at5r1O���T���\�'����ɟ���1��	�PR��(�)�e5����eAt�����B�K�D@����ʡ�_���qF*�HPZb�,Ѷ=��e���
��*�V��5���H:*m���"�U��ib��Z/C|Z��:t]c4B��AC��c4��Ɠ'O��^c���Y����x©P+���~_��E �;Ɣ��P@���,�d�Lj�$8��3�m��z��y������Mo�<x	UP����q�5NYhҩ�{�J'�ƣF��� �|{���G���h���_���M�5K�N���5�]&5u�L��;l7[)k����6��!�{���!$�6�9q�K�Fe+�}�<�NA�*�����r]�h����{�ˍ1��^]�IR�y�h�Vf���(]@����'��F>�"�(�~Gclnޜ,��$�PY���X�>֭���H�T��%G�FK���R�˚<�^x�P�L��F�H0����$@��-6�kl�lwl�[l�[X+��RR�$ݓ��d:��U*�hTU���s��S�>��!u]a�X��m��r�Ee��Fh�:q7��m���A��-��$M1
(8(��<!�b��1�r__�F���S}���PJ�$�ʹꘂ&�a<�ZJ���3ۑ�P��#��O�u=��h��{���5���[ū�5�,��o�owY!L\	5�hk�4�`�`��}�z}*�� ����5��56��xj�8?��ˋ�(>�4�'�!:P>���f�'�w��ƘB��Y�i@9 G �[��mh)[��F�+�w~Tn�-���")�"q�*�����P���Ze/��ѱ���f�Ze��/�*����Mq��Y�l�Z��A!�L�#$
%�)eB��ؐq�T    IDAT������ж��(
��"��O����L���7�X�Ob@	��!�����?!�"��h�|�2���}`�̜J^�AJ"���gğb�n����*Rʯ7�С���	Xn�4Е�I
( Зfݙ��y�l�;l���ߤ�߁���J�8g�5l�†����m�l���]�i���4E�:��]'l��j����>Ѩ�Ao�[���D�)0��.qu�2���0ͼ>6;y��}D
2���|3Mj�ZH�O���?i�@���3Yq �CY�gdG�,�g�2��X�<x<�M<���0q�f�\b�^g�h�=\�1�#�}oE5�넵��a���E�5��O.��9rB��~ˁ\�5��yX�x-��@QE���X�<�ji��!\_o�ǳgO�X,�Z�E��
ژ���_��m��?�Y��u��0|�缊�-���-��6�����粚�9�����\��p�������<�W�gT`*��]qrr�uAS��� D�6q���v���h��ݛE1���@�����2��9��rp���B�����18Ȍ���lquuc^�x�.�U��y�ꕸ��x��m�	�)>-^���3,�ivp���|Wf����R�\(���G�Z�A�8������k|�\�9��L�7C�b���J��!0�߉D�|���J$S�!����T|Y�a;[�sb|N��[���v�HC�'�!ZW0&�:�{U�=ڶ�v����������g���x��V�e�z�}�=�wX�N��?������/?�y��o'Y�M�˗��� �mՒL�ǥ�R�l�Q�>��������Jd��(�qxOv'$���|�3,��ӥ�L����r�#�a����.���%6�ЖV����K@����p�@���ޓs���u�*�E=ΘWWW���������h��/���Y4M��j���S���a��b��� 5O����i&�?ݼ1�ݢcw�� h�PDPI��X�;�D��!J�5�Xb�%{Xn�=��M��|&2Ї�,��O�����_��1�<�W ��:SնF�2���E�@ٔ���{`�e� m��}N�u��,͞��U�L��V�`����<&�_�Z�����@�yl�{�y������޽�_���ж;<{�ƈ=i�wx��Td	����\]]݌|Y��4(5IM�2ئ�Tb���+SI
 *:�)�
j�d����߷{��u��u��ŚȜ��[���~�e��J/g|���A������ʥ�4 >���E�����Mt�ezJK�A�)� ]�{��������SS���C6&)+�睎�SN��7�+C��xo��l{l�;��y����(%���u]���<j�����u]�b4�~?k��9���#H��_��)�\��.�G�P�R0Z����<R]+y(tG�Z�	�lc� AVeK��P��#�>
%}5�J��*�<_��M*6?����c@�5��EB#%��g�> Q�F���� lɀ���;[�����2��*���~#��t]��n�}{�-���Y�E���q������˗�t2܅�zkGg���K}���q�����$��tw��2�J�6�f�W��U�����J����B�<N[B.mڮ�u6��mo^�w�o|�rHr��S������,�펰ߟJ�Y��J��`m���m��_Ɉ�̄���~�6O�Z_�i㧌�Jz<�!0;��ri��ڸm<�7�W&�hZkU%���6����4����c%t�A�ǀ��԰>�J��Цj�s.r�J_�;
��»X���'�}��p~^���Vp���	������o�����w�����%�S��!���a�d%�~'�� u�qB�w��K�Fi<~}��6�d���a0��ui\eC0I�|�R�*��m������$�z0��ž��h5�~����Q���W\\�C۵��"o7K���&����)b	�*�������75c�/���!Pj�2�Ʈ_��T�&M��<�OT����gYD�Sx%��A�>�2ezHoˮ�}�o�,�#NM+q�<Bc���m���չd(q�HHn��B�r�Ç^�o�>ѽ*�(����Y�� R�f ^�@ ](��Z��XM�>X��'�%��@ZaK] ���4��D��+��z}y0�2[�����P]l%�`?�L�&�Q�t⇟X�r&���H`�D�g 2t}}��~�zQ�Dp9d�1���v �����#�0)��楛uH��^�ge�cm?��������g(�.z���;��-g	��6��Q��B�����
�{ImqE
�06���x�B����?�ࣀ�X�BaP�䴻z���
��T^K�9g#�`0���	@z��d�@��؉�B̚R��dlJ6���Ѳe����s��_���a(�kp����fW�T�hMZ�y*��d�I�P�ђj�!���m�c�`$!88��΋��_榒���)F�x�U����ո�!!%N"9�S�S乫��6��F$�%q�2{*=��Ϥ�%�A�ڱ`� �ǀ2�+O��eH����@�>�hr�� B�[�w�g���,%� $@��+��-Ҍ�Xs2^ěXGU����G����AA��MK�COcd�Ѧ+2��r,[��z������r�"y����a��ϟ�ʃg)sq&jV�@�@�>Q�OEB�1������<��m��TBi���
 %TnD&o`'&܊��\�q}=�gs��\�����3�c�(2��1U*��D�f�2CJk)M�'�d�>z��P��)���\�v�ä��T�@���%;�� ���8%�L0)��R�O��A���JJ��H�9kI$+�v��e#z����W���%�h�n��>��Ft[&0&��V��o�`4��6B�$�-Sy(�	��]�HUř[r,�^/t'=Џ[i��c]�Ҁ��bSix��fY�7���/�������P�"��i�c%��۳���v*7>{ A���.))�b���؏�}H�=Ȧ� ˥￾,��6����>���Fč�O:��`y_S�c@�1�� �:,ZG{MP�0h"�ΉO���4�J%���rNG��>��f�P��"�5d(��#5p�������C	Hi��=g�k�O�L�(���y��r(q,\>�n;N��sW28[��1���e�	���H�|ޫ|�%;���e>���y`��w@����ؽ����/���@q�c���|
(yF����Ӵ��r���:�$0�1�h,�9wy��1p�F���"F�JJ�2�t0�˜�=�ʃ���<�;���2Jb��TT<}���0�D�N�$���|]��(;'�ĥov��Ph��<�J�3zIQ76���}b�H�6���q/耵�X�|�M�!}��Z���M*�X�֑��3Ґv�Fe-�
^.�
�=I��$c�f.�Kw�2���Em)�@���-0A!�iy(�0ɇnxy��G�{�jz�1���V��F| $�k*�jbI����FN(P �c��A��0���bFh��R������g�<��P�
΋MJ��Q�� �=zk��ڮ)�	��>��Ii��H*}�	Q^+J�r��̀�Pf�RG)e�D�fѬ�(��<�!	9�`�I��PA�gmֽ�pS�8�~H�1��?�<o�|D�0<�Hψs�/�GR�c�J�k��97 'e09tf	|<�����VFWQO��6�)1���Z&ɡ$�(��\�5Q�N�	�y ��7FhS!�εyݐ"x+dR@�o[����F�3�����罋$8E�w�k	(>������Z�D��n���A��C"��nD�P����OI �$���f��P)�y}�FNswa�ҽEQ"����C������[�T��ɧ|ﲹ���i/�ݰb�#��7&�	�Rd�1��^n�	(��Fs!�I�ˈ�,琰���G	^��I�6 nUU+ �K���P�fN���f���$CI��8����?8;�	�_@�?���&��`�Fjl��y�y��ύ �2���y��A����L�S09�����.�4)k +Ys��!9�<K�*��Y��k��\*�s>��K|��_c@9h�3nk����A���|����vU����!��m�W��������xy�*�7����n�j�a���?+�.�V�(�9�|��6q.���R����,�T~���+�t��#ky�4�P�yMζ��U-Q"?��f�泓!u:#�2�� )̔]�ǯń
�,$���9I��(�jR0q�A+7gA�
��}	(��S1���ߧ�!�1�"V�l�'t@���A*ayΫ,��d;ɑr�զ�
�x�%z@`������P�	&��Q��:��&8��$�N>(��3d#_Q0):��Đ��BA�O�=O#�d��,�h�}�Q7$��)��c�ǚ��	�V�O�E �P(p�6d��#^���KG���Oʞće��8���`,h`}�a�~1z(�����A ݄��m�
�h7�n��ׇF��B@�/��֋�c^�j譥1�HR6��֢�-�i����@��+:�>�QJ+h-��*N.1A+]H��,��Z#�*d����uq:^)�"����4Lr�s��T�ܨ�����[�O���
p�p��KEb�[�q�2�^��N|q�Z�� ����	s��L
N��H�)u��b�)k��xd+%f�*S����Х��1$A&i�a�
�@E@a�*tmS@��Ai��hb@q��r��f#�5�x3�{FT�*�SЗV��C�JCi��)��6.m��8%�
����Ld��H���A�DHӨ�*wdT|��Pn������3�!C������:��Rׂ����p����D:cK��9��A��36�����\�Ф,�q?H�G#*#�0)mhe
�����3� �@0\�(��*Ļ�U�+�>�]���b�.��B2fUSC�!�Ɲ:���i�\6��������,�����ٕ�_���7{;���!;�e DD��9[�����<��o`�{GDR�BE����*�L�u��b�T��,3��L�T��"R��������m��P̷K>�� _�R��L��)�Q���T���h:<>� ˖���Y�>�8U)���]ަn�h�΢�A�b$b�|��)�NO��#�>)8����-��1�<@�-�'�7�@r���]��v븜�+%��a��Ұ^ ���y����m�l������c�DG�K��rn1[wp��=�C̚��IU�u��r����{�X붻����9�Z���}�o���m�F�*RU�MB���д
�E�U�4BjU�RChR��)mEr�H�
5H>�)D���R��P_>�u_ּ�K?�1�k������>z�YsHS���w�����������p֍�ۘΕֱ�%�teOɳkL�8[W5���RQ�=���|��sI��:o����=��q���&E�~�u���}Lo����k�+)�����nR"���0P����8]JtH,��Jc�Ř
�-Z��X[QUM�F���a��.a�����k?�0%�~Zk��a�Z�տ�W߽D(��p�zP�sVH9�ڮ3~zJDr���y0�2i�%E>x�	��s��M��9�Q1�$.�LMv�c� 畿�l��Ss/�4�$��D]$-Z{$S+[SU"7�(����ȁ
����|����\5kWq�Q�n*Sud��y�{> ��(_�}+*M�~5���qf\��o
��z!f5=?vi\�-@Il���j�Ȍ��m��P�z:�����SJb�J�ݘ�ʠ�O#�1R����
�<�${����;[D�C���j5j��gsL)��
ƔGkM]��Zs~qNS��_"��om/���,���A|f�q��zZ�YQ̼�s�����=��o�5�,���_5��n&�	������(VR�ӈ�+q�GQe:h��>�Ĳ24��miȰ�v�h��Q�GAG����Q ���������6��>)�����K��J���t��E@�̝ {%�`��.��_��ꥨ�� �7��2ˡK�JD��'^�����\%])Y�����Մ��H��j�-�}��������1�<���5��sP)PNwB��9�� �À1$���R��ʀz,̊��xb�����i"�%�2�1I�J�l��pΡ$Rنus̍�\�L~�g@��d�圣�;��ctv\*�>U��,Ɣd'��YiP�Z��})�������~�}/~g7������Ǣl���E]c������LJ�F���� �x�_�I�)�kGx1O��w�O�=:E$λQ�}¬�v� )��enn*�2���@��)�2	 ʼ��T���"h�L�X4�ƚ�U��h}ʍӛT�
���G@s��uݘ���V�2���#�9}?y[+~�G~��������ʊ�Zi��9\��c,��oL���	�k�d�氒��l o��U�]�6E��i`O�N�^�27 �(UT��}�ǻ�)0Y�(�6TUES�X�֬�'}���	}S��%�Xc�V���cc���Ik���6���y�W�{�./���|�?����������(_��$e�f�Fc��n��S��[�-T�kN�q�Z ��ݞgE!�+R�5�xf�[�oi��\��-��u�(S۸N�%:�1�$�Ԏi��[n��<Ϭ�7�TR���F)=iYg�ҹ)\��3'�[j��iۖ��a�w=^R!�h�X�fJvV�Dk��uc�Zl���m7l�6S�5ι��{۽?�����(_7P)����X������LĲ����\�D��\��`��
����.�nO�#�� $�i-y�W�tW�+iC���#�f�����o2��y�Hk=�m�tp	���#x������g��|����.��O)��w��l�`�A�b�Z����:�U�}����_w��_m!ac��l��	�e�1PyC��)��������=	Y��֑���ҙ��� ���4*�IRa������횜
I�R�E+C<�,�j֫��� ���2`x=�����nP,U�Mb�j��������%
�f�oL���P=#u6��W�F�6Yn^�m5�������E�f��n���5�X\�B	�����!�f��g0���Ut��)2E�d'*���ُ)Ɛ,i�Fk�|�T�)MȇR�LӴ��#���̤D�!��c��hͺ]�}�6���u��'�B3Iѵ\٣]��U]�^'@�l6��1������'�@�E(�1�u*vYk']�g<HW�'�|�%MzF`����j#������f"JP�5���d;!2ڙL��lM����(��, �U�F�C���J�t}���t�}?�J��R5��b�N��4#��=Y��� u���Hy1F��ep�n�b�^���m[.7�xҘ[7�7`������m��K��=��E*���HR[�mP��Ҕ�O���B�������1=�L�����'�?�#��1uUS�5uӤV�Hf��N��[Z$���r��,�,Լ jUeY��9>:�ٴ�(Q�������<>���v�Ѷm�wӦ�������~h�A�R��Z�
�~: S�2��T��h�gs�Ar$�CW��n����Џ,���_�~����?�4]ePM��� 	Np���5���<�K���n��,�X��	܂Y48\ޯ�V����>}�#gzfb��᫛��
}w1?طІ'gł�e��R,�G�V�&�*z0\Lk�\�W�J�K�ޔ>Nz�㤦�KDw`�Z53C�Ѯ�T3!������9忻���=7��{l>S��;���_ޞ[Pn�(�����g�1�앖�M�(&o³���:�b�5��.p��	\����b���wfJ�s5}��.�ny���n�f��F�Vv]ɼ�\��$_�?���<iWM:T����N�s�*��;�:=O}j���a�l`h���7cҮ78% ƞ�'I�xt�~0�z݁��#�B���>f�R:���o4ɻw�k��?��R�8/��f�->������?9ǟ���e��(��ad�oI_^3T������q�%�}\F7�N���x�o�
���uѴ�z]z	;Z��K�����f1�=�E��r����CqW)�Yז��D�q� �����;	�t�y�h��n�T�5�9��B��t�7"<��ü���fG?҄�Llt�p?&�j����>MQ=�dr�'���E`�<a�Nw��^{����Ok���6��ϫ���N�J7gó��8L���9���tԩ�:�
���%=�H
O�^��:���c���9�6�F|�}�1�?sۘ�@���k��dr�A<z�r�\x�8��v�w~�8v����A+l|*/u.��myV�5[\��,,h9K$��Kqy�sO=>(���;5h䪈I��zj�\��w���þ�/=����Ѽ+�䄜K��6���5���������ѵlm׶�v��8�/>} {z�����tY�47u��y_��O��8�D�-7X=�'��A������x��m��{0�rLɇ����=h22o�zc�4%1r�d�.�����!:��ќDG|?k�f�עC�О\^R5��[d47�����>ʂް`ړ�9��.S�fG��Qk�栄W���~����^�����Ƹ��L��9pˑ�ߔ2���eC�S>��������y?0ib�1���
�0�!,XMV
:O�1��+�-y]w$�\tT�.��umd��5�k�Y�EXh�)w�'��\���#�y�RN����������o�{24��:���w5�ݹ�ꥃ�[��؏�5v6��iIg��E=�{��r����!�H���0�����.M��r4E#0�����X���`���{�Gx�š�����q��W��3�)��vQ��R��[��ӻޥ-3���x�t�O�����c���g�숿��惵HNxor�S����5��.�5��V�-٪fUp(��ai��d,�zgq��5S��Gq��&d58��յ���E�����ae ���b��
�+v^�ѐ�F��>��TTb5�rDo�~~��$}�ճ�g�５��
4*8�C��U�v�z���=�ՍA�����$P��zuu���h��ʫ�%|é��S\�����п�����V�d�ʕ�*)N���3���tO�4.�[*�PKRow��+a�h��H��gB�!���J�������:�`�d��g	�J�`gw3L�K�9�䃾��Wm"Q�%k�X%PT�bj�"�g���G���<���e)�9 ����7��$ar}U,�1���{�s�/*pKf�w�G<ޅ�,!���꡽���z�4L��˹#]�(׫����"MV[&&*�t�\��rgSU�2h䘞e~�c"��Kbߍ=�ߓ��B����2E��eGE85�� ��8W﬒;��h �OU9h��ng	����Ě�'�T��̓�H�� ���4K5�ib*�	� �˩$�G�U�n�������nQ8qf7	PE�U@��:]_xD	GgX�|x��{���Yc�o�esYf�!rva3v8����@�c�]^FF&<�B�������,�p=VU��F��J��~ɛ���������Ǵ�K� A����D��]�� �������!./��b�&99�9
f�I�G��ʾ��vW��VZ�"+�f���ɢ%JPaF�ظ�l�'hQ,�4w�X�3�x��T�mR�+���),�Jh&O�)녲b�-nͬ]0�ہ-��1����(��T���¤�ôk��X�c���S�9]���:8Ke(ycB4@�/��o��D�
V�d4{�~H��Kgc-�ܚ'����fBb���	���e�J�h֩�t3o���Ș�l��,���v��b~i=U�����ӥ5���+=�3����9;iyj��f���-���6�n��`���߯�.%�*^�#=�Ĵ/�_é[��:t��[��~>� ?����?���hr�S��]�s��ݪ>t]-�.7!æ��?�i	D�|>���MK��hN�&�����n��6�ԁ�a<�j���9������C�ޠ�����{B�4%I�w$�Ŏ�2�h���L]ӸkR�'�%l�8bP���gi&Oo�Y�ӧ��Xz����Mf'�`�Q�'�:c"rx�%-��~�Sj�=����N�ɘ^<lf�-��6 t�����h�DU�@Ť��yx�uϭ����������h�x�ѫ�S�
K�vr�Q��
�������;�,�W���	��#�����e엣�g���͟��i�O\XtEXR 3���o[ۏHn(0�E��q^ʁ�YF�������q�����:��,r�ܘ��!��Y��$�OlX4<�IS)�&+�q��'0Hj	�*�E��1AHH~@�Ey�E� ��okgJ��a�T�)����j�+B�e_ɗ�Gl]��'lC�����/�ި�ߘZ���u�q��ТfI�	�#�Zw������U�j�k�^/ajEE��ح��N�ƙ��&z+������!�</mY�m'c&7C-��n�L������z.���=�6_M|�.4�ʓ�9;DR>+1ڤ��	��lJ��*���9���|��@	՜w��/�,%N�s���2�h��<c�RԺa�fǑf�+�Q�h��[��Hb����մ���CBD�#�0N
u%����̱S	�ǋ���j�1w�D$��[��8��:i.Y(˴"2x���xX�~�������#>u���?4�՞m��>W ����מ˨a1���ё���X���S�{x�ό�MLr�j�h�c�������m#q�{��������a[��v�˓&h%&.�Hu$���}.]6��~u;�����؏������O����,h��s�!��[�5���3�?95uwb#9�/��iF<
rZMl�'���1�׆���6�;h{Bp�u,e6+��eC��9��F����0�5�,��3p0�,����b۽�c����d rY��`|g�&fǾ,"��h0���ґ�8�[�OH���n_ߵh[ �9����;4C 	��h.���3@~��p�oc>�'��Ђ灅�$s�kL}A *�V����� B"�K��L#�Bݣ�*=�^Si-+��8�ǝ�!7n+>����n��Q�~sݹ¦�?���Y7�_
�H�-����n��������yY���B��pǎYt"�"kc�-l��t)��4/���#S�ay�\ڑ������iU���"��3!�ç��^6�@ ��>�(�}�
� ~��zЙqy���g��+�;�n��c"h^	(��$K�vKqS42P�.��SBՁ5QU�6qQ��%��2��<�#�;�\[�i�
!�T�D��T���6������n�z��Ԧ�����>��UV�Y��-*����y���A�RlZ׌e��IP�����Ɨ��92�;K�*�f篭�����`��}'s��!�g����]c��rr*���Lp�!�
�����qYp�u?���z�v��v�'Q�F#��	^�|��|1^z�hu"�I�ry�������i�ӫ��ze�.^�4ۦ�Jw�(,��4e�%�t:��`J��� �g'����e������C��GӖ%����3n��b2p�as�X��3��B�%�'g*����
n���2;�R�c~��[|�+��PD�fh�����m�C4��y���(��s��KJ����89p�{��s����{��I�B?�s��7��q���r��'�%�\V�e���W 7qD�C��V��5*W�u����9X��./���vq�I>?j�eg �_��I.\gɋ�a쩞��[�����o���o�%��Og�6�oG$��C8�7{[+�'�=9�9��d��C�P��>=�<nt�Q����=3+���<�nﲜs����N8Y����� ��dus:J\㉌��p���zfz�*zbe�3W��łB����='FG��w,~��%��7B��V!��CpC�N���<�I].I�b��.�h������Њ��bj4��I�F/��R����<3��\a�2�*b�X�A��6�㧀ty쿗�=Pɠ�#CiL��o4�d��I��\6�����=Oțc�m>n�}�Qj���&}>S��9�m�¢��؉Ο�q�W��u��_���?�xd��hoj��/�?JL
�=�_ξ�%��K�8}>o�[�W�o{�	ؼyb*|��t)ڳ#xrr?>>^��%��z�$�h��:~#�j��;�o@������V$Aj���,�m����f[�^��֖Jl.�C�)2|'�ӣ.�;Z��i��T���m��A�N���al��WvF�˸���b��9�� z�����[%[ww7ETS�|��,G��$by�f���Y<	$
��x��Z\��Wj���> ��=�������@S��,�O>�ul�.��^]	�ŭ����A�gbҞ��4>�s�:y��H�`?1��3eU=���h1�i̸�2U�N-1P������A���ݸl��y	�6��aY`���	��!/q�ի�������i{��~�~�n͕�w;cA)�ӿ���S4��`{�1ێ��I��U�Ǭ�Ǣ}F,��͇�pm�^ ��1��MDx�B�|���� &��03���������$�,YE������D�J�v�ٷ�ˎo����Uu�.�K:��τ�A{6�{�|W19ߔ^��@�#�}���"{*�QF�`*Q�|�}�ޞ\O��	�3����0��@[�c��(+��V\T�����7A����$�&�{����2����h��̽xZ�����3�0��6��������?������}@�k�v��F�)��C`����IIS�/�AgT/m���-��{w�娔���Qs��m�K���D#����/2��3?=�TJލ�nv�7���
�
>��.U�R�y��y�t{��{�p�X��?�X�ۄ�ߋx�
��nwљ���hZ�¼��m��ǯ��4͘^EEgA��1X������F������5�'�ͩ�i��ۑ�-*����
����@��>��Q��n�����U8�p���ș5�=ݹ�������C�Y�
����w���?Xa6��s����v�xU�����˳.��~d�Lߋ��]��zd"��M �m�^�K��9&<����Z4�x��#Á
����NH��}y�|^��	���Ն�<KDMr`��4�i�WǼ�פS�X%S?��5q��\>=\����w�#�>|�9~��w|��	D������m�-w�E���Fbt>��^]k�Tk�&,����逑�R��X_�cc{!П���~j/4L����;�8�?^��о�?~rѶ�z���2��1}��C��#�����O���zsJ�ݺ`�&�5Ko��?�)G�$�1#��E$dW�Ϡ��q��m���j|�֧8����d/���YF�5��TO���������pE�[t�P[f�"o�-�'�#����*?,�`\aY��Z��'^�&d��9H�k����BR��8}��_e�`���K�X!|�d�&��� � N$�@�u
��dX�4W}�B�DЈ0���sNRt~��KRq��8��	�[¬QK���q"�+�_!�I�;6�:�'mI���v��ґhc-�w�=x��(u"4.U�F��l�����*�6Λ��tp\�F�ir�*G�}࿹��k��V�~B�}�Iᚾ��N�^���%�N�A����;���U�AE��}2g
Wz5�c�5��<!�B�X8�xƤ�t�鍳��#G�
�3-����x��M���@ �����_^eBC�����B�8�"���#2k.���$L�z�1J:Ĩ45�v�PGK�D,|���8U%�|�׭E��L�;�$�	mN]@��~co���w8��;9��7n�c%u�_x�,R�.C���ϸGMK��oC>f8���W�1�ډ��jBij�*ry֖>]-�|��MVߨ�����s_���a!M��1���]�=r�k������pQɴv���\$��k���<!ݾ8�:2t]���2#{ۡ��\9c�0֜�a>~�UH=J���/b��᫔����Q^��������m˟��4��[��}���'���ADY��f��z�B��\��H�,�)��щo`�45��D7S�qq�g�*��S��KÝE�8�r��LK�� ��Q�1����$p���3o��*�h�2�g/h��#XQ!�{����|��YqF��6���dKC��L���6��2<IQ�
s\�Չ}���e��b;./֯է�է�p�� ��3p[|tP^��#=���1������{��{;���X���pg��C��8�d���[��,�� �3���>���N������c=�p`G_d���`-���H��i�C'�M]��嗏MG'���
M�K��q h�?��r/'Xv8��	8}��O��'��xl؎�
~'�/��d��U_��,"��	v�������W�`��7VR��P���[���~��z$2��S��>�%BO�^�Q���yQ�o������r��@t�:F��:����/s������	Ss����<�{�p�)��ѯW��u�J�ވ�م�T�3��TbB�Wij_O�GE��F����Xh�[��~o7B�鹴��~�5�������j��7-����hw5�ݥ�ޙ�����yo�nkf{���������Qփ��F��܌��o�~M{�D���Z����80�9�p���C��捜�rсܳ
��0���/�I���dZ��A� ��a=�ߪn���u����bK%j�TS�`1�L�m���{��uZG�o	��
��
+J�6��}*u�7hz9�؃���k,efZ/�P2�N�Fd���<�:�[Z+����I)#�dl\[�+=51c���sf"��-�����'�ఞ�@� �����`L\5�r��ڣt�g�f&��g=f�2�EMA�a{f%Om����RB[b�/�XP@Ŕ���O�Rx���up��I�ϕ��b'����"�}�-(x&��1=�c�I��K���A��/�\�#Ş�e�Y��r����dO��FV`۝U��f�z�W|".]v>9��̱
��i��%��ܢ+��qn���-�v�X�W�a��>̳�@Y)+�������d�⟚��������Ɩ�5��]p���9�SRI��բA]M΀Ž��
ccE��Gm~���S	�����O����:\�JQ�hk�𐆛8��,�h�`�Qw�K,��N�Un��S"��%`;i��x��㕃C��y�Q�����&�a��`���*!�f��p����b���s��v}dݾ/gz5�����[\%�*C0���<����{�(�$���@��i�k�x~�߄ZV�d�=<f���,�̠��s`/Qb�$gi��➔�7�*���]�z�C���-k�}�3k)��gqH���YtX����I7/׭Pk�.C [�B������G���8S����D��tQMs��� �0dE��u�a���SS�,�����ML��H a2� ;ua<sv�܃�\�PL`�=3z�$���~t@R���G��Y������ni	SG��@|џ4#`|�Sq��\��{p�{����%�UD�街U�%s���=��!�ĞN,Z����!����S0:�A.r�k�CЖR�r�w3(\��!u,���S��7��ex�Jy3�C3>�,'ªo��>ȹ����;�k&�B��"�;猊'�lu�am,���s��L2+��[	?~�#����Ǧz���*-z��Knø5��T[�͵�?0��Z��H��KM�QBa�_�װ<�EBA��\��B���L]�G3g�k<y�6,��~>ɀh?��x��)>�e�u�$�y�����u���|6m��1���Q��_�Z��7��S��Qlc��m���q�B��}r�6Ĥ��CF��ND��+	䂾`�6-77�u&n�E�@4����y��7����?[��m���� ��<�����ܑ��WM������7U�~>�L����w�蜘B�� ��F<��~�P�pſ�S"FW8��h�Qn����^Q���]
������[T^����O{�X��Y 4>�t>�����EV�jK��tRT�v	nȿ"M�[s��"3������h?1�M%���`�QkfK�1�׺���	�l�R�+U�]�p�t�dQ�����\�s\�_����I��z��+T>Tx�]gf��6�\'���Y�F;�\O
��^N$���*XN��:�x�s��(}�k�y�����V�_����i��֨/�>G�>�o啾�p�M?�̀���$��,11-��f� �Q�Y'�(�"���8�n5���ur��zR���O��Y���q�헾wz%�p�W1Q?xx'x�"LPU  �D>x�}H��%жL+��&uQ�8�w�9%���v����*G��� �q2�<N���L=�������c�%�������%R��}���,�>nG�E��N�<s��P!M�9 Z}FNɢ��n1��{˸j�;�	hOLբ���}�����ي��ZT�֙��,Ə:���F� �����!/%��Yxu,˝k�v��ƳT�"o�tݞ~�3�K.	�	PeV���R] 8�2�u�l]��A�s��T>Yi1ueؠ���"�������QR�gY�@����h�rm�G���{��iejY���0[���us��")9�im���͇�`:�Q�Q9ڮİ��p��U(�_���Ou&�&*Yga�eC�|�Si�s*(<P��&�_��J7�Ќ���l�]ٌ:�r����v�C�ߥ?�"��gL�8��t�E"�BQ���>2�6�)���.����z��z�m���b�5^�
Hb �IZ'��$���������w���lU�l���g5ГҢ]��`�0k�}�.;x�{�:�V��ɴ:�e���z	M��-��))���<�J�{/��E!Iؽ_0�� ��?�2 +r.��q��Q�S����gh5���euR~<,^�%W]�~0x��H�|��o���sJ��1$nyV��i�Dj��!�|�i��1��r
hƁ嫑Г.cvr�6�����.;��״����mXM�,X$ȂZK�˷�H~���%�D+(�¡V�@B	�X��V�)(bD�dk���4_���5�B�k�
�4����P�����6Y���������>?�@U�UD��F}&���������%��IE\4�-���HI��f#?�r2P�hPd�t���� �����K+�m�ꫨ#����i�q���8����61�� I�V�H_����pO�^:�a�ehr'Dm���#@���	��kc��M�&y*߉N��0qݨasK#�g�K!6*�A�v%~�F3��V|�+I�")��������>�����^�Y����;�"��B�u�['׹���c*�WF�N~�Q���9h�f��<e�p�ŝP����fq҂�Vwh��}���@�*�]SV�5]R^���-E$hۑf�����n�� /������k��k^~�܋
�������M�AS�Lz���Ʈhp9'Zk+`�A��k�����G��eǴ����3{�#?�Y��<�����t�C��	`�-q�^��xqFϪO�GDv���>��vt�B����}��̮�/Ӯ��/�Վ*l��a�@U�jR�l�T�$ƭCz���U�;�(ȼ�-����ǯ
�M�UQ��V^f��Q�g:��>�$���Qƀf�W���+��C2j��6�\p���J��I>�a���א� �}z���&��rU�+�4�LeF�uRt'�:Bf��cH�$��,�oK֏��q����Qq�i_[{5z�R>7������2��j�~�V��3�>����	�j۰��ϴ�O��(�e�Г�"O��J5�o�^�X.1x�c�'��w�t�Kk���*�3.����!�@�O<_���X8�_���U7�Pu���z�t����2��&���	Q��� �nF�$�`�Vk{�RQ:~�{Ķ��84�e^��O�{q� c����)w>Y�g2�ZI(v��rw��'��|(���@)�dk�;�Tc�������R
�E�,����F��^��EB�Dĵ�+o��i#n&���W[r:�G��`�Y��-�����2?��g0)#	�����7����$��c���2�hT׹BԎ��h�k�ҍ����K���Q�`p��!H��f̴�>2.������v��]���?w����SF��� cx�f�i:9H������Y.�1_�B���;�WȘ�V� ;\�:�mw��1t��N���~�﫸U=Y��E�H� _�Ƃ6�߰i*dx��*b����9�Q�J���p�N�[by��n���%b���,�C�ҭ/�k������Ȩ��S;���v�z(��鄧;e���ܜn�O!V��-��.�T�*��ц�rL33�H�e�Բ�-j}p�ff����)�lqQ�&���0������g��d�5��VkU3&��bJ9�Y�Ʒf	�B7�|��k�GŐ�03���@�Zh7�x�G9�zq�8�F�p�b�Bn�[��
��[�J���	��?��]R�ˀ�C�5ԓ��{E`������M�P��;^'Ŷb|:�U�	ȉy�P� �����Ұ�HV��b����W݀�A���ʯ�kM� }����&P�H580�vLY�%�o�:���oY^m諌-�j KO��;;��Z���bk��擴��3 1�XH����w��fEr�mM$��!<I 9���vZ�F%m���^HT��أ ��a�ÿx���n"A�$d�`0�wAǛ�[�}�Qy]���z62��g��y]��ơ���̲�����Jp�n���+uYyn�,7���a�GWCG"���g�wQ�{�&��¸4�s�f[�-�vrO*^���}sH�n�W��Yc|��⽔��ǣm!4�i/v㥙��D,�-�
�h�h�V�����w���qJ�*(x�&!YFVR�+��G���Xj�U�2j���N�K��"�$f���]�Qݦ?Ow��?г�(�4/�7��T:��%1~��Wo��Y���_�d^O��_�ƕ�_�ز�I�"z�ޏ)�(@����|W)6ՉKcw,1�w��K>x��s��2�z��Bvઃ`8����0��QP�&"�|��2�gIm�~�%e�����d��������WAy�U/��:�o��>�������D�AEb����@�uS�_P� )��Fi���Y5Okt�yn��MHJ����hd#'nl40�����c�� z�%^��,�������ʍ�a�7��ӭ�jy�1�d���+U@8ɷ��j��hydC�3( ��͈�,V���)�z�w����8i��95�*�lf��9�ZV��rcB��y�"�h?g|f�ɽ.�08�,iB��~.h��h����״��C�����is�k-�M�į4�����.�)�X������l_Ԓ��b���_y��sf9��c�LVi���e����#%���7v����FWu�DQO�i�p
JӷƟlfR�5�A.Я崺�����iL�ku��l�����֫�L��3��&y-�lG���O��"l�&;�1����.M�:�`��u��`���a9V]�_�Բ+Fr,7��C���dJ f�v�A�ɷF���Œ�KJ]�lޏ^���2�����˧�9����%�9y�Z-��?e?7�l��u׼�.b��x����q�$��2 ײ�\ִ&eȣLOa	W��V�z�-4M&X��.��|�L���뭎:�w�2� ��5oYDs�`7���=�[r.i)���M����0�4�K���bD��kV<��|�^c>2���cN�����N/�=m�c4G��^��!�)�#���r�S��?��3r�|��:��q��({*d@�'#����c"YKX�W�u��.�V3���jb�m��'=)#�Y;h��0������q*ط8i�
�� ��đ�1v�F叫�M�g���MyG��#͈�}CoH?�3H�G;���o!m*�_^뱭`hlGk�]�����o�"����bK�1U�F"'���Y�yt�g̜����U�U�<��H���u�	�m����P�[�Wi����'Z���Z"�y��$�?Ėe����L�'MiG�=�Ǜ�\}�c_�}N���/(b�>��:��\�~�At������ک���Ds��kK�_����@ϻz�(�wl$���˦��bN��?��M5P<�	�Y^i�����g�J>g����Dʥ��V��C[�d��p�k����q|ZA���f��W����YKA~�DJi�U͚9�7 kFU�ɑ��;)���M��grL���`&Dz�%��`�;�5l��
�]H��_6�=�ν�T�Xt�к��t���Q��= �� 0CÂ������a�%OxTI;Y<�g*�*��U|ϐ�$���ڌ0V`u��n�PD��K	$v20�FR���p���/��y�g�bqp�B�*U�p�@�;�EL�,�U��D��#|�I$5�C
� �x���R�WuY筛NV_A{NGG�F�9����3E��r5e�W͆'y�9�:�%X��Y�x|+`�i�y�mkj���1ykO~ x���U�V�-s��~P��u���|V$����/u��4�i��aS[����j��z(�/!7�����I��$S����V�ti�#4�'��4i!8�ԗ_�0UeI^��yWl�}�!5�2P�V�u����Jӯ��稜��V=V�����O��I�K��yM5pA�-ͻ��H-'�"��h�O.>�V���������Fd�4�lM҈���4�!i�'8¡�,�|�ut*�U]�����D��1 ���.F�oj#|]x��Y$����u����[(�?��S���(�7�0,`��=Q�nU��MN~ܴyJ������X@�F��?������F���w��7m�d�J�;�:,Ý���� Xa���N:e�����&��I�!�d!�<���-!N���ܢ�8�jBY�ʛL�P�#���4`
�712�df�����˚<���?�h	j�Kޚ��j�I�ǈ��)>ǹo����Y��3
�}��)�fw����<�c��&��C:Ho�y#��9�cTZ�޴/l���jDv&;��q��E%�6�;��ݏ�<.wb�,հev�nf�{E�����nkV�B>�~�Q߿���D�u;�؛Ȇ0�-�MY4��ٌ���I)��Z*f��\S�5q�x�q�̰~d��[�i��C2�w2��M����Z���Jd,ϴ�o�X�@)lo۟�<����>9��^��,�=֫�Ue�p�|��v���}?�3R����8A�~���)������o��z�y_Oٟ�w�5g3q���̄+����3�����B�Hc�ƹoʔ<RA��?��M���偮���u���^�YG��4���Vf�N-��e1�/��-ئBT�#��o�(T���(2V�͵�ϣ��s	`����)˷C�2����g�¼6�`���{B�9E�t�\#��޿�4��X��!뇗��ʀk]J�ߖ��f��B��b3c�t�=ɧ�t���N~��|��`E|�R�O>Z'
��"��s���<��CPH �m��K��C��E�#��I�s#�қ� �E%\��/�]`���h�_%ۙ��]��z���D�����P�v���Fs8i�Cė���-=�N�<<'���[�|��߫筂�C�țV���+?�Bk���f�WBΕWi	Ɉ��c����S��\M?'���(d3�
�7�0���E�Ò��6��1)�D��_����b&q��K��5��((�Myd�>�L^^c����B��}B��ي�_��^!'��﩯Ȇ"yAB�%�b��*&�S�z�,Oէأ{}�i�=M��Z��/\�(c'��Z�F�<!@u/[x�J +���DEJ, ޽t �"F��%������Q'��.]�}
X���ҷ��q���-9sy�F�<�� �|��`A4�-�H�`�O�q���`x܏w���Pӡi�$QQzsC�<�I��gP�{��'T��}� 1��@-���۾ز�y���H�s���;zp�B��R�Q:�t���bI3#�-�Y�{�a�����eP	0�xX{X,���2�X\�,�D���;.��d���q�>����=�ɺ��k`��Lu@�m)��ܦ��b\�pui�H}���G'�N�C<�?��7=�%�bf:��T��8d�A�N����ݫ�g�������o2�(�����<��1kD�*��<��52�����/�2�˘���UFl-l��a���w#� �[�_�1Ϣ��_�L���`�6��U	��_���?�#Qc���i��K7���ܲ��įc��R�v�L�ܠ���W1wIW[c�0�m4�8� ϷX��NTi��#���:`�C�2���/�'��|�f�,��j*)X܂:�J`��H���m��=��m��87��Ϋ�e�f&��͑Dh�U���h-������>��m�(��#R�}�4�b3N���9�b(����E��g��_�����ת�z+k���+5C���'u�*eI�o\͏-s�*�!�*x!����"�KG����ʥ����1h��~�u~����=9�\zcv�踤 ©��)r�pGs�*��@f��b�/�����~�)��f):ፘ��9�����q��)�ߍ�5�ˌ�����e��AEg�\W<5m������n
hФ���ӦE�$N�@�7u�)���+��a�>���z��	޿�3.����)��B-a�[�֍���v��_�[*{_�ɖ�Z�`(�BL^��7*o'���d�Y�+_n�R]oWzI�J���å�����C���$4�	��� �vŊw��	%\������[*��*��߯�-���wD.�v��w�o�*��힊��	ܕ�?un3���px�Rp��5������Hå�̇�� !����fn��[t]L�(U_�x}����	����cGs����v��be�7Ӡ{��)6��:�^p}-��hn���8H��ts��^�>��Lg���C4��H��������BZpV��sԔI�~_l�����v�����1.S��U��Y����P��Ee�_��n�yj"�Rʭ/��\�PB,AY�.�e{_��d�a��8�߸�� "S��;׈ƣM����ƌ
Z�GV�ڸ77kb���E���4�;��a��(�Ĭ�)=i�^RԀ�ؠ�4����-ЩF&�g�Dk��r<}c9�<���D�-˻WU�����~�Oix��]%b2�w���kgg[��a����sX_�� �w���8�g�[.�l
�LL(�ak��(���DTf�?�ҷ* �?ΛH����E�����a���0'��1�Iug6[S�pG�(�����
����磧rQO˨�mG��5A_����h]�N��uTx��^�[������۽���y�q�S����1���w�cm�S�hB��	�]�"��U;�"#qѪX'jc���u��@1�҃��]+��z��^U���tAS.�p؞lȏ"kDV���x�2����ς$d"�i8G�s����"���-=Zn�D�l�����l@���Uqr21~#�P��#�lOwC�ֿ��W����Z�WlM����r1� �w~��})�w6
"F���U�"��i1Ę-��	,a�g�6�%l�_��Yx��Ǝ|%�˃{��S+Q���:_1t���6g��Uk�<ɴ�:�Y��!�4�)����0Q��pc�\��#�.V����P�$6����-��Vo:7)�'e7tz�.�H4���F�ΰ�����P�c��{��d��CHrD2�Q�a�����^<�����D<O�:N%B�I��ܜ�(�1�y�E� ;9VO$Q�C$Mz��a8[8��=�[&���t�l~��Ob�R�R+h	Z���j1jU�ڛ�E�����B��*j�ڵ��Ԩ��oޟ�����;'׹��z=�s���gu�~�2�R��C�z���'��6��.��r�|����˒].l��r�CX�����]\�-�ށ�C����
4��}]s\?. >�QR�V��樂��"�=Wg�v ���p�%@b؅��MD Y���u����^�d;������.+*�f��ɋ�R�C���Ӌ(ݝ�e���0��/�y����ˠ�1:i=����Ό��qW��c�^D-Ų�,s[������/ـS�1�}X[�2`�����9+�}����,]'���M������yo��K.�if�Cy�����Ä��-,��(LJc��fEL�EeO�����nY�F[�
:�a�sḿ~v�D���s�'1	L��1�+�~������\����7�՛�����ZQbG}��5�_DjJue(}�ZM�!�K�7���;Y��|>��^����v����	e��"�u���|a(�T{�;��fY�f_3 ő`jL/` ]��9G�%ԕ��dd}�U^e������C����z�:���Y���OW�|�Q['dH�@��%S�af����W���W����NমqћI��u�~�w��յ��9�y+�������n��U�����ڎC���V柾5�^���^��v�=�+�����D��aja��\���9�^��Џ��>�Ս b��ER
e��}o��`7�;��9d?�G��׾�5��mM�ؖ��!~'�I�����٦v~�n�8}�ܓ�M�K/�7�^\C!1'Qq/�|򈃟<^$�`����3�����a��&� �b`#��a��,��@60ہ�I~� %�XF(?�p�?]#�P�'�ْ�}n�p�7��+�8E2��ж@�M��,=��lVz~��n��|)�u��<rG�EՃ�n�ǫS�m_0���T&���������|�*>k�Nz�8���h᧩Q�{�`��q2�9i�ʵ�̽77����Q�эk���lT���
p��#넗w���*t�1���Kgi�����S��@>u �Hʊ�Y<�Y\"O�h��3C|����]3��V�������y[M͑<mp�R��}�� �w�E��?�g���l��l7��C���Y�ǉn2ʑ|`�τ���������F#
x����Bb��p�C��w	q�g)���`�+���:��]h�|[��R��Z�eLH������ZI�)5%�#X���[������Y��J��vG�*|~ٱ��;1{������W�!F�ſ�
h�	ং��Q�@���W����	���HL�C��V�Y��D�6���,'CX/���'��=I;<��]����oz/�y��0��kP��A\���A��U�zۻ�~a�2�� xϼ�;�q�?k��>�3c������:©��,A��L��T��p�Ԋ��bs~��T�P��! ��C�*z�
B�ǽ��s���Z��>��A8B��!G��<�d#�L�l��zAn쐅&���_eN��� �׿��Kg��g����.�W/�vh.nODv���r��S�Vh�j����I�Ť�n�R��P`�Ul����I�?����Y�Ͼ�`e���uC��#T6~�A���6W�������Qd���md�i]��a��bq������<��\��������m叨v>�s����a��r�_�0N�����~!F�y}���ᴭ��Z�Wf<��^�G�C�zy���uT��	��VL�
���R��M5����*�f����X[�/s�bR�!�OM��u�

�t�3}���C?،����	��O�~Pfm�4�%�t�ɢG�~��Xa*���܈Z�ۓ*�v�G	�=�'���Z���s1�F���|�����|\��A�2"�)���gu���:�_#B������M(d�3N����7sG��t�0��>Ư�����m�w?`�w7������l@���Z�qt�-���@�oK#�Pz������j�`�P���|q���%�i�2�ER�����×*�^���,�Ol��j�c�����#��ц��h�s��j�qa�r���a���`�|I���t7����T���#�W���OU_�����V*$6���p��_|ȋ,�n.��;s���MA�p��GY�Р8����#���Wp�����g��[H�+\!�&��b�E�WA��A$L���7
�gnw�l�޲��� �|h���aT��<�e�x ��t�H������4������?��}u��MƑ������Y��>>EA�:{����lй����
3�c�?�7��y�c��T��Qu��]��`�v�7����n����?+���oNʿ�z��2:���2�T$�Ë.v$/�V�v�U�Qt�ޭ�������W�׆�:?�OɄ�
��O���Q����o��<�`����M`��HBt��ghh��#��������QU�`1��O�%]H>�����e�l, �9����}筯{��46���<�:L̍i�d��������M$�����ع�mkҔ�Y�[C����ٚ?G�� �C�V��Qc.�JGW��x!���c�����ߟ�W��Í4���SmS��)�	�cW3��3ɺ��'�g��5�
�g�6\��B~�6q���Z�h�6h��S�?Tmӯ�# 9�X>z�?�����ww���T~�����
$�	��q]�}�6���/=�nN�����F���P������h>�<��,F3�_���$��q������^�1�P��$-0����Q$�YR��+�Pst�o���_��2�n�pӑ�8S�̓�����jhw��_�k5?�*������@U��_e��H?v�S���}"�������e�*�I�"鰘
	A�5!��,��ۢ�)k�/�Y�]��ɶ�o���M27^���?���\Ӭ����'}��`3:������$װ�!���:���¤:���������?2#VXew^��C�P�ܩ����p�^��C�0Q��h�v,��h <���2�&O^�Z���pj� ]�h��qx���vd?w�!ʞ8�)��[�]"��4o�q*⵰	���b����r���ϷGo��*��=|Cn�a����z�%蛍��K� �c�&T^�c��yt��5[�)�P��>�+S$Q�rҁ'r���L��GXU(,���}V��%�<�"���.l"4�"|b��	/�[��~�N�����iS}�M��z�h~%D7���`O=�`�o���$�� �6�ʗ;U��QjĹ��yi�ВceY�ڦ"d�ZI��6+Y�=Ԟ	�P^=�ڢ�ږ�N6�F��G�Հ=y��ch��@fz۠Vp��	9.�KS�
w���ԑٽ���Bˆ�Ȇ����VqrXRF$����ъ����(K��Y���Ll��w8�`~�l{��(&�}r�!Q��2�S=����|`����_���D���� �0G�t$�:��-K�`���AP�C���2��V�h?��_q�t-�xW���3�B\r(`�#C���Q� �j��=���-�	��3�>>�iר���{3�Q�(ps���d�l�Љ�5�B,(7V#�
�0]�/O��|�W�C�9m@��d3�3�jCf\���l��\*��	i�%��9>7�%0ރ���r�2ϫ+M���Җ��Gx�b�S�����:I�".�c�yԚ(٢�w&[�$��������%%�y0��}�S�������,a���p�L爥ڝT�w��Vlp�&Rm�D/�j	</gΝ��c
=�9�XY�C'�������m.i*-�!�x��F��T�*�A>"�J!W|�z�)����2�Е�k2�MÛ��!���T�3{{}|f�0�ѩ��>`O;*�ݿ�#�msV���4,`�V�x�f�ɹ?F�W���AZ*ɧ�i��k�[�؀>�Y�������C�CH^��X2�J��3�c	�V�O>T�je�q����6���^���ބ�U�R�<a��%-�CD�6�"��v���Y2�m�d��\\��˖��f2�8�Á1�8l��x���7�X?�g��H~߾��O�hv�c�����>�:�s]A�V�����Ł����̆���a�1�.ۭ[C��W��ؔ�?ݎ�Pr7�q��{�,��w��*i���G(�B�( !�$�-��~I+gZ�m�2ho�ͩ��⬢p���xɕ��s<}vR��u�W���K�l���xJr;�B�K� j�<����&3���X���嫷aSQ�&բ�����'~bp����	��Wg0�E�R\>�G������.7:��Wj,��"�!C�׿ߋ�*��&�ȼ+&F��Y�D�Ȱ�{+~�ԖuΑ�op��m��D<�g��RNͿ�i�k��Ǝ�t���H�hi�"V?���y��y�{������k�C (��hqqL�c/)E�:��F`3x9m���}�`�q
WT�7�5�+%�Ni�;��H����̿�u�&m�L1�.:��e.9�;c���,���n^`���+�e)�`+�k��e��G<�k����Zg�B���@q5
���x�@e\{Zb�e.��8jJiJ��d��CH*��׷���dz�a�H! �ylE`��b3�1�[V$��BX���9�%_9>���:Hȅ5���Ae�-Եp��3{�"�vr���{�){��l�����mȒV�G��>�=g4T����ӆ:d���?�J�F[A�~����D��2B���AkG�b�����yf)8�Uv��(
�&���pndN����y.m�J�-���t�+���$-�[e����k	��b5>�f�h���y�1	�Y ?a+P���1X$-��s@��7?�ؽT�Z��"����w��tqt���l;�(f	 �Sĺ���*n�i3pS��ꧢ��/0����'��2 �2��.���Q!"���+z����jb����m���E��0d����4������J����]�/p><��P|�G��ԣ���dW���:���j�� 3y
�$-����}#l��_<6��- �Z��@�Ǎ���xXn-�N�T'K�z�z)������nꮔ��d�e$'ȷ����(����{�o�	*���W�LH2~v[(��f�q8L/<��4�2���w�>��}B.2x�!��
|嚹}��ݍ�Ϡ��Ͽ`VCx�w�i�E2�1wÄ(u��z���-�ތB���ͭ��r�ʼ� �hO����$}�G	�;�/��Pò�0�%=9��$�Pt0t�l�ka`��p�p����`�ly��TUu�d�N,���4���Q�9[,�G�5�xk�B��0��7t�6���U��7�'���Т5J#&�A��7I!��Y��Z}�w�.�'Ŀ��S�>��}0�u|j*�LD俧p�����(PM#߶��a�.M5;�0���q�iV6�[�l����ywF��ǧb0�T׉���l��kB����c���l/�:@���$C��DS�peԃ���piI?��f��u�p5�KУX�{#v����N�| �ٶ^����>�\0���M��Z���J$y���xH;:��Ej�GHx�3�H!������0_�nT0�)�p�_�g���~u�[�ؼ�eJB�N�NSE7Bf9�Ē��ؒe{}GH/�Sd���o��E�f׬j�8�|S��R��	
g��}��`^���w}.��噴T7���V
�?�.�%qXn�맚1'�L1=��]I	V�ɀ�ίĩ�?��N����=#���X����e��5vq�ycש??4,�Fr�t|��`;<�R������h���H���u0���s����xv�G�tXb�(�N���gTߔ+v���SP�j��=�R�B�R� Z�*��+�@�aWcS�e ��S���	�6�@�,����n�P���v�ђA��p�t��v�~��}4g��8�-I�\K��T�2\��K�K���Y���U����Q0t�l|��Ҫ(y�#[b�fiV�iN��q�9�p����j�K T�&��p��F�;[j��;&�[ -h�y�#�V�������e��X�[?�Q�u
�IS��t����㦳}04�p:ڞ�n񚂯��4�g�5'F��!P����}9B`*��џ���٨Q�	CG�B���H>����er���̈/p�F�cyNm���"#�i�K@��6��\� D�S~i?�;E�W��C���BD�h*�t���x����V�U�g����iU43~EM�l=� po�����E��� �r��k֮q�k�A���K��ᷖsf[����Zn���Ն����[Q|�+��'����-A�� -������YC�������;�yN�!�'S����T�LͯU�> ��(���?.�I�Xl{T�u�+R��Қ�C�,��I"�����Pj��`'�������t����+�P�Ǥ���-�X�6?u�a�͡�S��e`�RC��$�B hN�~���6ɰZ��6���ۄ sk`bA��.�+s
��]�Yb�x"Ŝ2�8�r&At����~�Y��v	fA����XCc"�w觅V$K-5B@������8L��\������=x��aV_3Yԓ�|��ç�}~lq(�j�L�tq>�:Ȥ,��S98���*��!B�Z���	�v QL�q[�c <skf!w�<*����i߈����'�� »9��98ݕ��}&6I,�Rr�U��W���kR�u�}����}XZ���	�'![�6���p����3@3bڒLٔ�OW�9uvp�4b�hA��vδ��G������T���⇤F2r�j:�޷p��I	N/4.�K/�Ϟ:ET��
�y��@��<���fy¨�n�2߸$\+�������j\�)�+�>��+��E6x�[sSl���D�}�Xw��t�I�WVV�`�
�2=s}�ta꿠�;��x�[B(?4��;�y�a9�9n��.׀&39|��@�v��ݯ/���H�n��r��A+���m��|�o��KW$�3#;F�'��\��#Et~��H h����Ltޢ,�vB��� m8~vA�	OR�Va�B���aL�!��H��݉�U����0]�&�N2|g@8��O�w������TrO����8�*�����o��=�ښo8j���sO�~̯�X�!�9D�3 �]`�#����(8p0S�����C �~�$&s0/mH�ǻ��Z,Z-H���Y��x��o]j!�ykI�����m�T{#c!h.�v=R���:R��O3�������C�$uc��g.����J�Q����:�̓����*6�?�)�`�Z٢ߓ����i"f��n�W�L�/3��6�`d�ӥMӱ�c^~^����l���b��Ӄǯ�tXeY�%��Nf6S�a���,|�o}���A��ӹ��v��l� g�&⓯߯<5�^�V�ϟ�㯖i���Ay7E����2��LDV^��5AD>�iL��D���1�D�޽Z����щk��RQ�cSܗZ�?�f����}��8(��U]/�5y��h��F�4LH�*�(��ͻ�C�_J]qu��DE#�0���2�~�İ�O�'��śⷾD�U>Cn$���C��@�I~&:։�I�y�\�������%�b�󛰅�@�'r�7�lP>�>�>5^�q��#�r|\]y�tN��$vE)�/�H�f���(d����s�hZ���=1�@�_�?�q�}Iۯ��ʠ���dU�"0��!ZJz��H1�!�:�b=���C��uE�D�h`=���qpܘdxu�"9x��<N�p��{鋈_���o�ӣ0*� y<=e鄠gA�@�>pޘ�"poj �q�-c�Ә�F�v9b+���EI�:S�~�����[s��T�o�AK����ů���p�Iw=t��oܴ�k��2n�(�'F�G�F��T���
$�1��%�{��/Ǵ���_�,~����&�~q���|b�����</�-�Wٗ��-�y�$h����O����B��t�Q���*l�KzFc�I!.o����H׉a��[�-u���s��'��6��Re�������s�.�h��\���&����w���N%�Kԇ�jh�g?XQ^!^2
��0w7c~_q�3O�D�${g�>@�4�H�Kc��q�c\�5B�����^��k��v=��/�_�\������Ph5��T���fy�ȼYn�r����vZ#�S'�9+#z��eszN�P�� �,�w�2kH�g���R�m�6��pG�����N>ΐZM��&��K5��UQ��K�k(~�ի���Ȇ��lS.�`t.+���VV@c�
RиI������՗i���Wo�[2:-�O��-f'R�y!D�(�"��ȿ�#�CF3�J��o��F�U���J�2�3�P�j�k/��aM��\���=����ſK���:����|u0� b�d)��6���6��{��� ��s�x��R��{Ǡ�� ��y�އK����qd5�Z��g�t��?,��;^�-�H^v<v_���q�4��z��Ⱥ!����Cz(���<A�j�g�.9�m�e��c���Ɂ����.\�3"��Ă�?j���7L��_�F���J�L��R�,gGo�R�.�@�v�3>�`yNeQc3�b!�	���fN��f�ѱD�-��#�LԜ��|r�ە;X�گ��E�M�ш�|�w,u�Bh7����G�i���q��ֶS�����X��dqG�;�hc���'��q��n���q`n�^2G�5+2�dV�j�C�D�8�sq�{��/#gq�#,dO턠�g��V)$u�5�ck�e������u���~��RT�D�KA�):/(Sey�R����iগ�ǃ�3�?ܱ�X?Ι�ɮ^���L���F���5էQ�H;�����Q+y%>B��w�ՙ�����U֏�����#�� P�qxQ�gם�F�QɡA�FZ�e�F&w����Hu�ӧφ'��2�������܈,�A;�gM;l$/��B_<I�NWQ���z�L���X��Q}yƂ����eه�9/� #bRX�V��ljC�CQ�t!o�?�C����3˜C��:ɮ��(�2����n���Z���su�J`�vݙ�m����]�������K�ǽN�'�M��5�9xh��ݣ�N�@������L�����?��-L���\���AV�����?�ry�Y�� �Ԁ�l�f��uo�Gi|j!ˎa6��{y��bM/�&�5*
��������9aP�EY�@�F��Aʁ��O�GN���w5Di���x1�SCH�b҄Xՙ��,O�<�7X���(&wX���ı�#�.纺ǂL^''[�{ዟ9���C{;M9@1������"�9e*�����m[*�3T:x�`Z)|鑝"�Q���Ķ�7���9cs82U�wއ��j^1Z���m��3����O�{Q2�7z��?�v��U~�����G�p�Q#��QC���Ӡ��gCC��b�bb��X�6D��i,�9�{����� ԉ� U ����H����&L^����o��*�A�B��P��y!�P:R&���mzR�x����K>�w0��P�j���5�`���G��b�ս �n�Q��Rŧ�IQFg:/�� bR��k����K�/6O�b灛>D��<�eF�6�S� f��ŝcǧ�OX��8e���[対>���}�����(	`<�4�6.��B�	�r�?���f�\	�`�3�V^0���0��Lݖ��l~�k��q���<�pAy�2�_O���^��V"�'<�	.��1���IԲc_�i�8W�X�ښë����(�Cߩ�;���`�i�+��_���?TnlgtK�D�ÞF������g�,�X�V���@,@ ���)c�4��%��5@e"�@|�����P����	�� '���ѺUYmׯ�_KVi�n��b���~��	H����CHq�OI�xuM^�3Ȏ�C�հ��_�ᚼ�7��}���ڏ��"ds8C��r��C]��Oً�S	�pU�������5ȫ�1a!le�A\!B�8��g�����ʅ���I �#F@�'_��Lg��4R�t��I�������;ّ]Y#9�5	@�1w���z_+�m��]!M9�RLc����	gM���amAJ�k����O\O�K�Y ���C{�`c�m�<Q���~Ȗp��TT��(zȜ&�o��i�Rm\Oyw �e'q�ؽ�9[e�/p�?��!��R���N�-���CϽ>���7<�X�\�H� �(ٳ�7���o=�q&�|����j�:s�����&���E.<EJ����s�Fq�Z.+B@�Kj)m��T� �k��Q�O1���j��vƢl�;�:
����*����C�� �k�"3%�1�
�_��4�3�`�̟O������k�&�?��Ӌi����3J��k�W��?~&��*���-�-=r�o��h��ߎ��C3��m��8ŧc�A��j,3U�x6Jq뭢ذdS�Ob�v���/��R�,����ن�9SO��i�zU���`)�_+�>�>U%�v}�B�cjJ�LC�Q�@fև��F�$ �Z��H��;�`:Wz��v������jqK����Ԃ�F�}��*��71r�w~�qz�T�����pN@��^�. I���I��8��j�ie�����H���@>id(iP\$�c����.��E�l�}�k�G;о�c�Q����n}�|�ɮ���� `��|�kx4O��7=��LT���-�K6��2N��P3�JJB|2���z#�t��Q]X*�7��J��︥�2��M���荭I��G8a����w�+�>�j���|yM�������d����` �;�t�Eiu�������1�F���Q��h?�	�\ʹ��6�O8�b����Gf��aĖ`��*�ؙ�.�%}�ڠh�Qa�Y?c(h��߼7���G^^Cn\NH�J�ת5�]���i������Ph�oA�	�z4�{�7/?�U&��<F���.�v�U{����鬣�H44v�)f�=��>�_ŭ7.�=��q�����E��n�+�h�����0���m9��6<����1$"NKg3�o3����$%���Um��(Ȑ��'�$��r<.k�����z?�+`��c�N��,�`�$д!�7`YV�+?XY�J[|��\�.+��
g�k�-@�_��N��wlJL�/�^�}��]ui��Y�5X���FM�� oϢ;��W��{D�~�:����h�EzV������v��a��?�ɏU�CS|f�^���v���Q�=s��5şHyH}V���M6��߳�f9xVw�T�4P/�	Z�v�՝qh�`@
#��n���#��S��Ǟ-����WIoi(�ɀ5s
��y�����/~c�n֧����|�9GїOM�IKB��V�ۭQ�=����.��꨷�cݯ(d���&).<N��SaY�N���F�����5�-�K��!���i���� �wb���t��v��a6>a�3��1�'E�S4U��p�x����+ ۡ����Ώ���W|㴮����]`�n=QKeA�����B�F5q�O	J[���C������B��'����\nF<H+��ץ���d�=:?���q9Q�*#E;��,�nN��'�[���S�5�sɎ:�������ҿ�GM����N�Z����o5$C��8���w��,���.���̊��,[�a��|�����zI��s�.ɜ�Ϟ8`W��ş�g���xV({~%��Ukt_/��P��:P9��3���ju__}�ɍ@X�MO]��,2T/��!h��|�#~��l�bQ�C�z�����f>�37� aB\d)��0M�rV�u>7�;�}�R�p�
:�^3�������K�;�����B]����m��D�D�:	Me�uA"O󧈆wB�5���e�֝��t�z'�v���-).%���7~�x�s�ؑ��o���O80�<{�R(KHh��-W�8�Eʁ��qG4��>Jb���~Ir�j=i/������N��M�O����I?
ŀ���:VN�#�t?�>Е^��ȫ�3J��R�8�*��|���` k�����cVz��λ�����窎�>� 1>6ML��F���R���DJ.��(�۪��F:��}�T�}�6鼽֝����[�"!����ao,R�C*�<�2!7�I9�L�^)� ���T��?�r�)K2o��9v̏��}㩯K���z��A>Q������	>����2�ut�Ip��|�[}+$�I��!���T�9�}�y=u��<լS@#|
���kj� 7�w�j��d-����Lf���^��
 ����^&��\S	����j�G���a�{΂Xn�?���('�b����	T��U��W�<�k���U8��r�(�թ���o�O�(Xу������x��6[�GT��/|�e����R�OHe�K�!|��;\��.>�i-4Z�VHԊ��h�YqVVK�Q�idH��.�0��@�i%��k(PzkY�ۛh��Q!�]���uɥ������M��gXsGc�P����y>
ن���A{ѓ~���_d>�%�����ց�_�A���Py� |� ����&n�n�uf��%m��un��K�:���"|rbׅ^�Vl�d��`�Zz�Ky�8##�����̤� ˾i��AK�?�<����a����S������l�K�	3��x	u�+T���;�����	�#$��t	�=R� |����g���Uz�����:��*��G���f��ȅd����d�yDx0;5��Q+JyG�3�{�Z r"�8��1������ݭ�mmff��h�m\X��{ѳ�pgaz�oӭ���F��e��ʳ�uLY�^��6���ɝ�׏u�Y,�*�9�>	3�z]0021�˗�*�$:Y0��m|��� w:2�� �F]�̉XV���*6|j����z��1���&i��fo��,~�%C8B|�n��aq�F�*�*���<*S��DB��ɕ��lsR��4>韶nBr?���R8��v��¾��Tڶ�Nίg�#P��s~��A��FC�|A���z�k���־��Zr�By�T,��
���y�A�BN@���iϨ(f��&�L2�}Y���h��*Q���U˯��Н����Ї��\>8���)V�ݨe/a�Q@�.�īo�f�}�_l<~��(���$�^���9FP����#t~,]���Y뢮U���ɓ(�2ѯa8C:}��*��`H��Gg4�X��[i��OLdFR�2�?��ZLM�J?b����[��x�Zv�U���$;1:�����Z%��cf�[i����t�i�C������
<C�ۨ���ǧG��,����3R�jPdI�^מ��)��]�B-q:�ԏ�7�ႈН��̓�4�&���z:�+C�Q��?����V���i�r�O^�J���΅�?ĩ��{L�����WK��i8<E[�L�Ս�����d���$ǩ�a�8!��\+�xq�f�f��l[Ў�q�7�v��y�����X��45'=h]�9D8_4�m�ʎ�ܝ	�6��g�sJ��|�M����m�Sk�^|d��K0٬2���\=������HX�F�o�Y��>*2�	�<쫢��U�]"��ƌ_<yw�$J����h�Џ}��Y�c��z
vΒV��~�quRs|Ƅ��V��v
w�p���>�Z2f;Ǚ�6��&䴲��ϻ��bw.�G�ms}��u\��47�R��Ԁ#�.��1�8]��T�;�m$m��40~c6[�:�œ�c���������u�z³����J����╰]b�@Z��� m\�g"�t+?L�cގu�2" /f�3��*��� ֞p����<GGE��S3\x=�ɟK^�|\$�^����*��覝��� ��'8tD��W�4)�Nd@\����e������a֑AYDDH����s����#�06��g�����,}
;���v76�{�w\(4���w243�������0p|��{�q�|*�u1(��W�y�',A��������H>*6�_�yF���*}�x�t�z4�w7�S��~�_>��nۓ�'��Q��/Y�� yF�<�2q��$�Ă
�L�G!Ƞ�ƺ[��c�4#�]a	SZ�'Z�e���&�$�1^��*�x�/Jv3ra��amr���r��3������<�ߠR�`~����b.5
�DO�C��0ns�퍠&4��$-�xo%�"�l�:m��������r�Oak�o�흊/N�Gb��*%�.:fY����;�>9zr�s_���8
mK�����^o��6q}P�.ŠΙz�^ajF8�Y����O��{��Q0y��AQrN{�l�w�˪�1^W�x�_�>-��5�<k�M��fN1��z%��u�������D?���}RB*OdF�C�ھ��r�=Z>��@��-�ԯ�.����˼�gK<Bj��W'�^[��x��Xw*�Cˁg0�tCab�����>/�Zw}A~C�o������t�nC�"Oβ�tw?"!�Lۯ�۾�B���j��!Ir��0i�0���y:�K�}���?�O�y3�����l!ze�^Z��'��$�$��mLQ�o��z�b��T���2lT�$�C
@�r�e���&xnxȤ��c(��P���6� v��s�.�lG��r��!���В ��Õ���ød�;+h�@��M��XN)Я�Һx'����$�|Xs�[�.��EU���7v���8� ��Bl 9u�Õ���MN�Z+��������
�l={��E��8��5�����Ǘli�ӿ'�t"�{�X���������]Ʒ�@犦��E1ə���#C/CM��(���(1���{�Y�f�K�3чWV�X=x.]u_�dM)=Tb�J�zA0r~���b�"	&��v�����D4X�ȅ��8�M�����5Ċ��/�:��ʪ�wC�������Q�!^�N���Q�~�����&��o][giD����OD�,�i)�W��V�I�ym�-��(��SP~���H8F?]�󑵬뮖6�!��w9;��F0mє�����fٜ�x[�c�!�j7�I���ʾ4���`��صy��B]��*��(Ua��q�yTV/�n;M��<b����/�x�7.�O�>k�2�b�|��ؠ���j�$��?��<�{Lm��!��b�7�u¼���@S��B��InEorn��eƄ�9�|cK�-v؏�f���������߿�����~Vu�\E!����s�X!�t}��u2���݋lA�AZ�@���JY+���`���N	���xf���z���d�*h�zsG�Ȣc���Q��2Q#���3a���Sa�l�+\S&���l�̸��vj�3�g`fQ�;�Q�U~K�"00�N��ۛ�b+Um`?y]i�� \~s<�ܼ�x��#�Op���S������ȫ ��@�1/�3|�}=�P 3�/.9�Yj��k(2G�E����ٜz�S�.+���1�4�bA?���jJ����w�ͳ %��>�Cl�R/��Diq_.6yݿ���+�uw��.^^����oމf�b&B	�`��X�:)���Exl�N�'� 4�räs�2Hn&��
6�t��t���$K��~��W��3��$wku���o	�^^����qę-�Z30]9Ւ��'0Tʗ�hsQL��s��=�+L�2��%t��>�8�J3&ۅ��Ѳ@D,�,�a%7���c�JI������[G�����8�y���G^ʗ?���Vo�W�Z����v��#�{�T��&N֎s�fԸ}�kuu��z'�.�C�٩�v愃d�^�>�"���a���o�AI��:=�~4]x�y���y�q��p�Fo����"�X�����S�3
�Woic�A��������ˎ���>��#��K�%j��v��ܯ6Ih��ٟػ]õ�ؓ巗gRL���g.R:.oW���̡�r�����ը�j�B	����YZ�B*��4Xϵ�L������e{�q�u�=�Dń`����~>�Z�A�����ӻp��}��8H���6�;`��wҸ�@�  ��z.O�:¥��Ϙ����KuQv7�z��~�ޏM�+������5�D�&�h���B���pM,Q��a��QESA��k�o����s�G�v��s{�vy�����qNO�9���4���(,V��uW�J�v���\�f�vW���/����q$�������������c�HX�opw?V�e�i((�S��
�_��H�o���I|�������L�VUN�^j��MU������R��������9�������o��%Qa�N�%6{Y�Un�0|xvYr����o���'��?r��w}����ֿ���?پ�����X�d��&���|�x��g[uE����rϷ;�n�G��=�?�*o>��{l�G~�����ț��7�lʕ�:�����j?��x�����|��o�����z��ϓ�/��r�<���#�ڒ�cn�]_�7��6v���.���������=��ő���U����<�-gԔ.�Β|K4��#C����3�8��X�]�i.e����]�P������W�xj�u��������Y?��-����6T�3
��t�d�?�<]�\�9%4 PK   R�?X@�G��  �  /   images/e086d210-4fa0-4a6d-a74c-91bedc336751.png�5�PNG

   IHDR   d   S   i��A   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  WIDATx��]	x��~gKf&�%� � ���ejdq�"j�kq� ��j��
^T��P�u��^�EY�"��JI !{&��������0YH0�@��|�Lf�m����|_� �0t�h3���=Y_���i���m�M#��4�s������U4nF���!��V =�id9�1-�E��4��V�v3�c�C¼mEy��K"�� B�e���q�F��y<h���&�^�����z:$}d���|�zH! |��� <4g�z%��]"���3<5x^$S���@"��)@��%��S8jw�0ә�:�N�g������A�;�V[3�d��y�K+Rd��C���1�'FF1É�N�e��p:�p�{���AP�=yU:�d2!66��8�t�(>���s耈)2a 8�KJ���q���{޹�((ܑ����jH�����ג��<�n�͂Qc� ��ض��r(Q�L ~�vi��� �_݂���X���I��TTԨ��P]������t�י蛒���geC�y<}ߖ�o��j�f���_��˳?C����`�Y�1OLFj�I�ϢE8���z�^�,4��H 	;H{FF���qǽwchE�wCb[x��R]��N�ҽ��=
C�>�iv:��
ґ#g�톾W/$̛���/+�m�&�j��38Ll_HQ!'+����~���ݿF��_�UR�ڗV&��+��F-qa���}Q S�d	�G��}�(y�(G�g�PQn������`��X���(%fDGG����Ɵ^���� ��u3�޵�L�-����ia�a�Iމ??�>�?'��,�fsOx��A�@�,�y�i���?Ěի�mhM0B�H������w���Сx�S'�7m��ڠ�~�z����cѫ��dF_}��J:��ڒ��6���>�����K �icO�'D,��۶���������W���m�gk�hHd���G��u�t8^���T|�\b'!�k�{�	,�?���F#"��f3v�����t���An��( ���w݅Xb�c��po�M��#P��K�NEjvVā���%&{�{c��p��G�����A@x&��1�>��I�ᣇc�,��	i�={��� ��J�Ŷc�`Է�'�TbP�J*��+�������0E��	6��+���u�\����d��s�o���&?����~؁�(�QT\H���v5��pbF���_�ݷ�p��~ۭ��yFD�N�};�>��Q�5h�9X��1��B2��C�;�h�˫#`����P@��l�	3)�+k1��7�#�	�3%/�r�ˍ	���c���o��˵32���I�{c�;�#�ԟ�,D�mE����ws�u�ĽU>�iRՠ�h�~2���(N��c2 �#�S~��A� �f0��֨6�\�����ܤc������Q}���j��A
�
��:�r��^?(ҷ#��o��ǩttPC-�*��o ����,D�MC���X�J�_�.��OR$���O��j�E�i3圤@�-����qaQ輌��p(:� �|=̥q�F/3u�|����+S0b�>�H��>��ŀ��`0��$�{óyKX{* �x#�,-q�"1�=�U� 2i�@#hͲ���o$PF�v����	yea����<rq������A\��2�������]`�b5�A���k������'N"Ǒɠ#@H��'0�Ĝ�#���%X�ȗ�y��!a�'Ӷ���'���3�q���1�sv���P��t{��	$F������������7���w�|*�gA��W�X�#F�|߽���*h��ڭ�{ֈ�-���i�r`<d�8p�̷w�N��j���XS��R cL����Q4>�7!`0V	)0W��%}i��*T���-����JD� ee���������
��jU��i)� �q���m�/���遇�6����oh|ri�9�F�rs\R����k)�E%RGUU����b1����E�]��눝:��>��c/K�S��b���~BxPz��n�4>��N�"��a~�)��`)��m����9{�@b���jԯ��aW�t�DQ��ó�k�<�0*f�
��r��'-N����s��^+�wZw�f�	< �H!.�}���:��	���X�<�
�q}r
ي]�~�Q��dk�6 v���#��S��MG(�DV��,.<��ޙ'��uW$)"S� �����ͫ��B�e���u�Lx�l��&$ f�x�-Y*`��d23=��)��M�F`�J��p��vy�����O.��U�H�(����קk`_�������L8��v�т�	�_���Yk�^/�1�Eۦ��X���"-�q�g����Z�w{�
9=Zn���M�0q*E����t��Y��TR�>~1D��/L�g�V�n�ѣF�|���_u��pD9�|�$� ��<k�"�=��dۜ�p�Z�G���p=DVD|Q��Q�"��C|~N��\W�,/���F�ZA�%���T��c���-2�] =�%j��Tř�6�/�9����E��[��^Ty:(Hi�P[V.y*����s}�t�2�a��6xSS�����^�C*�1Btj=�-�ȱ'���W�K���6(���/*n\�8T�hu����k74&3��E({�)X_���T��B#sX
q1Ы��=4^�q�ƅ4��$y�+6�#Rp��}�/@�����
$%%A����$��D�O�X�v'��{��ߧ��Q�)=k�!i\O�,p���Ʒʰ�nv�t��M	��0 ���ge�WJɐy�Jv���%�z���E�2�W.�(Z��r导�RTM=d~#H��}��0���]���C((��ك��ރ.6;rJ�;$j����S�&�[��S�ݡ����Ǩ3!t"��N=�&I�
�8����"~�$\���E��i;\`h��zŬٰL����+�^��X@�a��h�l��'K|%j�C�X�hx� S�z����'�����С�f׮Zk�_Ҩ�[�����~� �Y����፞��ER�D���z� �
�s�h���3���e|َ�Qwm؀��݊ď?Fz�y���e����>��Ha8W�Ud~5F��ڸ�I�ds�ə'�1,��!f������`w�b�h�p>+9�,���"�'!��7bI�Gkמ׀�%�V���Wk���9%�S=�a��ٛ#R��/�ƛ�E��u}u��^��C�g�ҝ٧KG�Č8p��͸��[�զM� 7O{>�.W8j��UxL�7��������Ld�w��zH�D(2�y�Å^
���-yb��^L�c�Jt{�=\7jV�[������	T���6W�z�ݱ�W��k�g��CD.��8T :�F=�	�.D�|j=D۰�����o�z�z�=�J��ɖ��G�h6ׄt�k�hh;Q�׵k�����ɬ�I���|J �u�ӳ��yB�W�Y�������3n�,]�.=.?���������C��8 �Ν�u��41�'��
2�����Y����&?�bz��*К/2���g}�]4d�*3ޗ�!:,��1{���F�+QQ�u�5z��bO�3:���77rN䬣bi`M��"�5�rqI=��̎��coT�� ���>����C�SO�|�T҉'(�Νa#�˧τ�{"�X��0@޴}�z�O0�	S��8=`���b�~��D<H f��/�{�K��gB�r/8�nraoH�\Y�=wC߻�h+�3 #!,�7d��jT̙);Z�E,m��	��'
h����G���u��K��W�ܵ�8�|�!�b7�'&��J��A��>^���3QN��>B7�db曭VL��`'ƕ5��@���y�;K	�d�ss ���Я� G��[(��ӢNR���l��t�Ĥ����c�<�n�/p�)�&�Na/��&T���P��䫑0n������Ͻ�Ο}*��E�'�"
�(�.X�jN�E��g{a 0'�{�7��cͰ{���q�����cas#�sf��B��a�^~������]�Q$z�K.�L~��y�-������(7�4�w�/)�s�{�{m1�[��&���|��K3_|�eK��B��e(%P._�.��6o,Z�*0�$��%���LF��Ͼ��'Vs�u��n]�K��;�}��Q��vڟ����rY�*|s`��у�:k� Bk2����8>γi3���2�s^l�2�	��R�I�!*fÖ-Ōy���($�	��ǻ�o�D�<x��p���p���D�I�K?����X��UB�iԾ1K:vL��������U:q�� �W����\��rɛ���" nJ�hT���B]���/��	D��?�Ao�����7IR���(m���N&F=RT���r�b�h��;�nim|���^�@�2�_�~qd�;��"e�=�g��Ū*D/i��KK��$v� ��w��P��)���@�H��<�(I�O�l4�Ȓ��"N�{?��8�	��}�fa�mu�����>q�]i{ϒ
���ݞ�j�R`,1 �8F��;����&�xK�<}9�^�W�~�g��� ������@��3�0h�`���4M7s���0�"��Ñ��(�4g"�t�^$�;�C-�R!O�虩���N<�ܳ�b���b������@h��e��
�D��L��?.E��ݽ��c����x�z�tf�3�B��]Ϟ��j1��"UՐ����!d�G�j�;"��:����E�"~xu5�yyj���lWH5T�^9O��$�[H}}���ȑ#��
g#ƒ���x?�������#�{�m��&H��[zZ�<R}π��B�ˮ���p��O�:x�P_4��G�č9��<\s���kx0B��s�Y<k6��.�z�!� `voނ��-áh�Yl i��h��Mh�!�����$���w�����;.������Ȇ5��>|s�6|s\��cF��8^�a
�M�!�7�'$�oN.����U�q�%��h7������A�؝潸�dP�(,���ųm�s��x��_�x�H��QV�(�8"iC�DC"�w<Gl�d��ۓ<5kb"��@�F
���N �LZr�ɶ��~b0x��J�8v�3E����!�۫�YY%/��0����P@b��F졐�'��L�Nu�RU48"���>��덐�s�R�2�\�vȹJ�Du a�� �s� ��\���5i�ö�v��<���N���HmpS����M��ƨ� "v� .[��E����Ⱥ��xi7�I>�ۇ� �:��mv����J���u��oqڀW�j���I`tP�i,Z ȿXSMqF��    IEND�B`�PK   Q�?XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   R�?X�Ti  F     jsons/user_defined.jsonŘmO�:ǿJ��u���黎�+���B��8ݐ�<1�w�'i;6wކ� ױ>=9��>�����kl�9�Y^�4�_l��U	p�C=M��C�`����Ù���.���jvyv�n�MU?���47ue������up=Z��Yd�h�<ȡP�&�c��I�Ҙ&H%z���ӗ8V�1u�i�A���|�8M)bFƈ�$FJ�Ii#k8F�pS����>�	z��K���
l��̪`����*o6�~<����5y鿨�~����RW��DT����a9Hg?�j�>�Ӽ����?țein����� 5�Nl?���r}�
���X2��i�.�{�����{'����{a�:�l����,dWN*S�U��b�T^���/+C�?���b/����j�^�%v2�1ӡ��L�.����_�/�:���%sCǒ�~���n�XPԯ����)���B�G��	EaO�j��Nh��a��6@2��~�Cb%ca�]��5��X��ġ%|�n�҉C+�ź�:qhIOl�N�Yʓ��ԱƆ]ۇ*�Ա�(�Fn�Xb�a�Cu�2t��b�T��H'.�IuˋN]�V�8�"O�[\l��T���p����y��g�W���D,�Qd���3������IF56)c������|gv~��
w譇�۔���E78
�G}��wkw����<��6�"��U��Ia������.�}z\+�˴i���wKo��,940�*m�^���,������5/4��F�[;����Ǻj�u�734���4/sh��~���n�7��/�ʃ>+��(ΐ�8C*�©&�)pX�kL���YL!D!j�A<�V��i#EFDb�M�ep�NE!�iL����R����$PD|N	XX!"q�`<��t������~G��+D�R��P�Pe��m$�X���ԑ�:J��ܠ�$65�ER�]1���>�E;{��b�~�[s�JJ��l���txl��X#����4(��2"#Kb�aKtE�����%�T�,�h�����S���H��e,��(�e�%���ԈqjOd��O �XY����I�vX�,�H2�ZB�H�Ư!T�J��D��*&��4K�~�Y/�^?_?�PK
   R�?X�O�:5  �.                  cirkitFile.jsonPK
   �?X-Q�� �� /             b  images/2f436d2a-342e-4b79-b795-89e98e9450c4.pngPK
   R�?XeX�^Q3 P /             3� images/a8051118-2cec-4f18-9b89-ac75f15be4ed.pngPK
   Q�?X$7h�!  �!  /             �( images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   �?XLe�� b� /             K images/d88fff2f-2870-420d-8277-ad43f3d18502.pngPK
   R�?X@�G��  �  /             � images/e086d210-4fa0-4a6d-a74c-91bedc336751.pngPK
   Q�?XP��/�  ǽ  /             * images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   R�?X�Ti  F               l� jsons/user_defined.jsonPK      �  
�   