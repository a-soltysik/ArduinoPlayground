PK   �>X�
7 �  /    cirkitFile.json���ȕ�_e� �D�n�H��/�,6��$�����ȱ��ԫV�g�����3m]����n��9�`�1f<�"�>�x(֭O�c�c��6�cS��ow���J���}}�~���-7�}u:T?����O�sr���I�Ǧޮq�JҶ\5y���$�2$뭸�^�+��*�۲r�[\�y�|���\%f����������`UpU03X\���
���VW��VWf���J3�U!�({�4KD
@���J�K�D���K�D��L�D���L�D��M�D�Тw/�9|�9���
���r�$�+�$d!M�"s���]��7�M勅��k�؋n'q/ps���c����P������s�o~0��J�{�[�{����
2�+���o��0KD
�������?;�����a�p:6���o��0KD
�)�Y��g���~����f������f�Ha��f�Ha��f�H�La����v�%"��v�%"��v�%"��v�%"��v�%"��v�%\��,)��,)��,)��,) y�3�k�Y"R�k�Y"R�k�Y"R�k�Y"R�k�Y�U��v�%"��v�%"��v�%"��v�%"��v�%"�+2{����,)��,)��,)��,��^;���^;���^;�����7�[��~7`�,�`�\�z'X�t��s��z��A�K��]��J'X��!���wP:���s�w�;(�`��=ֻ��N�t�Za�[a���	��Uֻ��N�t�*�ޕ�t/�iDV�Q�W&�Wf<��,����^P��d��&�l"�p"�t��0����P�|��;����S
�O�|z�3�?pR��	�O���N+X>��}�`����'`��w�C���Ew)�'�ؗ'^��.p�h<0���tB ��68�`�̧������O�|:������+�����Ń��O�|:y�8�`�̧�n�����O�|:a�8�`�̧S������O�|:I��K,���tz�?p���	�O'Ɓ��,���tJ�?p���	�O'#���,���t%�?�^�;���#��?�|�ө�`����'`>�t��?�|����`����'`>����?�|��)�`����'`>�\��/���O�|:-�8`�̧������O�|ڊ �8`�̧M���'��g���G � �X>�i�
�����0��� ��X>�i������0��9��X>�i��8`�̧�e�����O�|��8`�̧�|�����O�|ڈ�8`�̧-����'��g���G�8`�̧m������O�|�p�8`�̧�������O�|���_�X>�i{6�����0�6���X>y�ofk���s;s�v?��7s��&�3w?�>:s��3w?��9s��F�3w?�9s��֘s��u���`ѵ��G�`������`q��yl�j���XP�#y�"��fʃ����oʃ՛��o�݊I�{�h=2���Ƨ������2�+�ʄo<x�������.sI��uҶI��i�J��ƭ�~��g���g�ȝ����ۦ��pA��z�%��6��O�,+���:���k_�M�ن���-���6)�r�Hp��9�7���'�>��m�EVI��=C�m��̷I���^��i�O��)�w����_W��G���_�����B���"������1D �n�rH�[�C��0�����1D �n}sH�[�C��>������A%W�qeV�V�QJ��� &X�X�F)�멃�`�[`�ԯ���U��`5\`E�W�����`d�R}�V#���/շ���xb	��V�QJ��� &X��:�R�W31�긇�q�R��9�	V�=�T�ԯ�b���{��8J�_!�au<��q�R�z:�	w%w)V�SXG)�묃�`u<��q�R�;�	V�SXG)�볃�`u<��8J�_����V�QJ��� &�5q�EqX�:�R�W�1��x��q�R�:<�	V��������A_���x��(�~Uy��g�:�R�W�1���}�	���������AL�:���8J�_����9�����5�AL�:�������m���U�U��
�����@_�g�``�
��V���}e�
��V���}e�
��V���}e�
��V���}e�
��U� �@_�Bau�y� �*�W�PX]u�; �
���*�G����w�t��|�r��p�p�V8��Ѻ�HoI���8�K8�K8ɋB+Z�ל�-'}Qh�C���s��$0
�ph�����F���a�x�IbZ���\���4F���)�x;L9��@��K�8�LIG8�¡�9>�/8��B+Z�����(�¡�9WoI߈����2��e���(�¡�9po9��B+Z�����(�¡�9�o9��B+Z�[���(�¡�9�o9ߔQh�C�s]9�rr�V8�:g�sc'�Qh�C�s�9�rr�V8�:���-'�Qh�C�s�9ޒ�V$ݮ��e)'���\F�����x��eZ��j����\F���J�x��eZ��j����\F�����x��eZ��j�����(�¡�^"o9��B+Z����(�¡��.o9��B+Z�Q��4��4����'�N.��
�V{q���2
�ph���[N.��
�V{8q���2
�ph��[N.��
�V{jQ��8��B+Z����(�¡�go9��B+Z�����(�¡՞so9��B+Z������惓�2N.�8��B+Z�e���(�¡՞�o9��B+Z�-���(�¡��osN.��
�V{}r���2
�ph�g)�[N.���4ڙK��t���2қv�2���>�3UF:o�T�=Se���L��~�3UF:H�T��<wԁ/f�-�:W3~ǖV�+��c�Ε�����\� [�sn�Ì��3��`F��*�se0���� �WN�+�e�/
;WS��E�K�Ε��ⱥ��<?���2�$8_'!m��h�&��oܪ��	g5ST0,�PST�=�ڴ^.H�Y��$��&��i�eE���B܄��I*�����v�!)}[F�m��i�M$�z���?�2I�Y���"�$M�@��MR��6�Ґ��24�v�/ST�|�d�ӡ�=էfq��^v��ʷo�N���!��@B�{�"���3H�u�,�$�T!	�.!A�@B�K["����$�!	�.QB�@B�O����ڸ���+�(%ׇp�v�x��\y ���+�(%�_��0�j���8J���T0L�:�au����=&��7�V�=����\M���V�QJ��چa��q��(%�_�0�긇�q���Pb�8����:�R��>0&ܕܥXOau��=X`L�:���8JI{~��`u<��q�����1��x��q���4�1��x��q��Ρ�1ᮉ�.���x��q���u�1��x��q��έ�1��x��q����}�������t� �	V�3XG)�\5��M�כ�:���8JI���`u<��q���a�1��x��(%�3c���V�ǔ��̯A��� �Ba
��skЪ@_�Bau�`^Z�+�U(���:@�}e�
�5�.���6�Ba��A_- 0X���Q(��@`�
��U��hU��V���j�� �
���*VWz�U��2X�ª�s�'qQh�C��6s�%�.R���.�/�$/
�ph�^s����E���3���(�¡�{�9�rR�V8�:���-'�Qh�C�s18�r��V8�:���-'�Qh�C�sc8�rR�V8�:Ǉ��'�Qh�C�s�8�rr�V8�:��-�1�Wb�\�9��sr�V8�:��-'�Qh�C�s�8�rr�V8�:'��-'�Qh�C�s+9�rr�V8�:G��-'�Qh�C�s]9�rr�V8�:g�sc'�Qh�C�s�9�rr�V8�:���-'�Qh�C�s�9ޒ�V$ݮ��e)'���\F�����x��eZ��j����\F���J�x��eZ��j����\F�����x��eZ��j�����(�¡�^"o9��B+Z����(�¡��.o9��B+Z�Q��4��4����'�N.��
�V{q���2
�ph���[N.��
�V{8q���2
�ph��[N.��
�V{jQ��8��B+Z����(�¡�go9��B+Z�����(�¡՞so9��B+Z������惓�2N.�8��B+Z�e���(�¡՞�o9��B+Z�-���(�¡��osN.��
�V{}r���2
�ph�g)�[N.���4ڙ뜏t���2қv�
���>�3UF:o�T�=Se���L��~�3UF:H�T��<wԁ/f�-�:W3~ǖV�+��c�Ε���eB��`F��b�se@53��V��+��ckAΕ�����`F�غ�s?u1�xl��2��u�K�����MR4M�xWJ�7nU�����)*���)*�OmZ�$٬�Y�n���4ɲ"��|!n���$�g}Y�M�ن���-�ʶMʴ�&\�q��M�g���,K[�u��U��Q ��&)�|�di��u�v;ŗ)*Y>/���t�6��ñ�mZ\����ݱ��n��M��v��p�6��՛7����U�M!�Mл�KQZ���t듛�>7>}i{�����T����<�@8���Ť���t����/�α�p�1<�~{�8z��������*/��� �� ( �N�.,����Q���xZ��;}����S}j���/?ڶ��N��n�]\}��=��,M��;}2R�%\w�n�0K��t�Ha�p�EP#�Y�uQ�f	�]�5R�%\w�Ha�p�E`#�Y�u��f	�_���-D�D�O@�@�k��:��PCPD����o� �QR���Kp��#��
��vg/͙��@�)ŷ���+5��j��b���̱r j��b���N�r j��b���вr j����5\����pf���v��g���z��]C��8W� �4�S���p �i
��vmi� ��PO��*	���PO�ڂ���PO������ފ��
��PO��^���PO�ڶ���PO�� �� ��f�zj��i� @=� �Ԯ�ӗ�o�_a�i��v�B
� ��PO�:5���9���5t��POs@=j̿�d0���#3�	�O�|�Lu��A���	��U��8=�X>�j�J���'`��7����_/�O�|���ߠ���b�������_/�O�|��v��A���	��U��-8=�X>�n�F��|g��������z���#�$`BA��h��JбDйD��L(hB�M�!:��	M����=D0��	��d���&4��Z��T���&������
�PЄ��c<���n�� 3�:��0��&4�N@_�F�0��	uf�Ctl
�Pge�=���B[<:�xtl
�Pgà=D�0��	u&�Ctl
�Pg!�=D�0��	u�Ctl
�Pg�=D�&4��\C{��)`BA�;��"�&4��D{��)`BA�lG���&4���D{��~�:��蜒�s
�PЄ:C�!:��	M��{��s
�PЄ:3�!:��	M�����s
�PЄ:#�!:��	M����tN
�Pg�=D�0��	�� �CtN
�P; �=D�0��	�{�C�<�DtN	��9L(hB횁��S���&Ԏh�9L(hB�V���S���&�N+h�9L(hB��0C�0��	���CtN
�P��=D�0��	���CtN
�P�"�=D�0��	���C��z��ztN��9%C�0��	���CtN
�P���=D�0��	���CtN
�P���=��9L(hB����S���&Ԯwh�9L(��\�q�q�����.�n��1u���N�3�t(��������Ag�?��9w���up�+`��%��
XG�p�����>�Yh��u\W�[��s�(�\��.C5W�:0����Z�l�B�O/�6W�Z>����Ģg��%��
<5l��2�$8_'!m��h�&��oܪ��'�(��o}����)�?qдi�.\�d�^gI��Mj��$ˊ�'�'Ϩ&����_�M�ن���-���6)�r�Hp�F�M�z�I�?��m�EVI��]C�m��̷I���^��i�O��)����y���o�յã�.>e/��,�ц�Z ����.Q��uU�"�[�6݆��覢ۊn,�����*�;���u�i�^���=���u�{x�#�=��.bL�C����s�c�a���h�)�σ�{t׿5���L�2��'W�����Hw��dH(��,_���]�D�D���D��(��nH�g��L'���S�ө���͵�ca���A�A�=$Ç�������C���塠Ŵ�����۷��zw{R'������|�k�_�U��V�M{�J�)��9���OZ)?u���x�i��]�}F|���_�nFnO��^��}�A�G����;��7jV����~i��n�>~������j���&>x����ݭ����;6�y�;6���)bG�?����ޜ���)���= 9n�v��$��nw��!��&�x����e��^��Y��]T�h�u\���8�W�m���uR����U�
A���w�/��{&Y.����oz�I���ḋ*uO���Q��qs�|y��8�-��Ľ[�G2?�Hz�����}ȍ�%��^��+�+H���^��N��}��}R/���ʇG�b�=��|9��_Ž����r9{K/o�s��ۥ2m;����I1M�� ��]�S�������������v��wq��H���pX7{�Չ��N:�mw��eh!��W.~�Y?���ߋ���u�~kVQ��>#���o^w?�?5�N�d���9D�L��L�+������O�M<�6�]'��M�y��E�v�nV�:k�Z�}RLIES>)Ώ�r����ĥ��#�Ń){��������v/��7��ި�e{��w��`y���P�]N�2D���������w�����޸e��J��g!����y����'"o��D�[�e�ַ�F߽�.G��ݯ�+���~�����ݯ�����Y���n��|�~��oo��;���#Ȱ̖���??��X�J�
	e���2��UH3�Y��iK+�,˓u]���*F�:K�x��jSl�zұ4�B���ԝ^_<��e���[�2��=z(�s��C�g'�%eXO��u>�����:�4x�+��!��q��4�����h\O��:u\���u���q�Wuw��#���"�Y��ύ�E
��ww��{U�?~����C����/:���G��-@�y�l_���ݱ9�~�ˮ�����F⧷����������WR��y�.�o�)u}<}���n�=d��	6��9�%�N�X�ӳ����:����]�_���s��O�է�����o�.��߷�w����hs���z���N��O���er�n���Y��7{����s6��@�v�#��^�b��΀��wM��y�_;�-�&�*�����fy92�K6[�iƹ��=`J��ɉ�D��e&�6`���uݶ��;�[���b��oq�����U����f�{x�fS̄���BO"�Y�/c�6\��;|p�\^�ll\�b�G��f#� z�������}}j��2�lQ����j����w���Çߝ�����}^|�_PK   �>Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   �>X�]��N � /   images/907530ff-a8af-4c9a-ad67-f4101e76dea0.png\�<���?�m7vk���Flڭf�e�!�]�m5���J%���ӧ�P�l��˖��\"�k%��E����0Hc�����������*3����y��9�׸q����/v~!$$��_�)BB�K�����l��t�5}�>��;-_A"�E��?��Ղ*$$������iS��7�g�M��{��y9	�h4ŋn.T�sN��^��xZ;���:���i�������`�RaGo������oޭ=&�����O��)�ʓc#ʓo4B���&�*��.���C�7l�|�돯��b�z����+��^��kY����зR�k�f��IB��>&"↼y�G1Y-nG�W�m����)����}CVܔ�������I�
;nX��r����K��}��	VYN#����� ���V/��)k���rG��]c6���h��S�T}�CV�)Ly����Z�li�Y_��ū��n^���LL�JH��t�3�h�=+gfR�g�n��k�^^*�0�K�����W2R.hɘ�,3�8�K_ZY�&_,cqO��mW�!'(2�:,I�1:嵆�����^��S��I�������[���^�]�Sq��K&��$M'�IVi-��ۧ��)Z�w��C���w��7����o���>��~�z<���h[[�aZ�z�7��0��.�6������AW�x�z+#U�v��\��ڵ�iܲlzk��Vobbb�J��������$jp��0v����K\Y�+7n��S�1�4{;��1�r̒{�Ai���o��z��U&��Kq�,�<O9�򱪴���Ɡ�x��_7A�������TU��s�k<Ե����)��Gs�)�p�l��U����_{1�58�
;�譓���y�>ۈ�j|�MjBB���i<j���Qe>,�6�h����dУ�mh��E�Q�����Uޕm�S�#Jb�U�����ըL���賫��2����O�h�M<b���%MtW>�njjڣ��#��	���.�A?/�P�o�(��(׻�����Ǡ����?��*����Kݣ4�4í��)����I߈��6�^#�߾}k��QW��X��4����H��9�FwN��~m�%7*i���4��e��5i�X���]_����G7v�L�����JP9T�1�s%���b��A:�k�\�HR�]J�~���X�,�<`n�]vG0��+놴�x~}��D7x8[<����=ޔ�D6�0�#�f�?;$����*]LMMYѻ4!�d����E�_�e��-lmul�	'H�
�7��F��}d�+4B��U>=���]�>�o]48�\kK�kva���zյt�7�&�0�!���ۢfôs�^����)]|zk������I�*�<L$K6��|w�מ���<��F�ݍ��()5��ώ̽�x����g�2�27���a&w��LG��a��N��p�ܪ:�Ru�)��Hw;\��I��%_��8���8�hڳb�A�>R���4w-**jϋ���S)��\�O����)T�3D=��#����d���t8�Ӝ*[�g�SZ_��������b����7��z�Z�o˾�/�gxv<��ܵ�^"99�����Ѻԃ�0!F��&�k�����m�K��{�L��߸��V�).ٹq�S�TaG�m.��͍��=���R!6�{-��%�f�Ҋp�tAs�%x�oZ�N�-��N2����ݻ`W�"~�������N��E%WV��N�$�D����ip\H��0-�����,u��/[f}�ڂ�[J�2�!A9e'�	&$mi�zK����p��Ǳ�3���B� ���r���F=%��ꐠ�����\=�������9x�o[ )���tE��Ǐ�,M���МL{�JǏo����Pg��f�'`��6�٤��mMH6ゥ89�Ǳ6)΅]����������{���x�<6@ou�s�����԰{��V������~�*ی+ X!��ge�?t�޽����.�i�� �{1_P���ޞ��s����.�?�z3"���7��,��# �6�GBh�1�,!��<�UU��7�����W'�+�5�4�q�$1�ꗖ�4c#���&K��s��<�
O����e�l�����G�·�?+��t)�a��FżO��31�2�w)�Gk[�?~~}J��)��\\\Ģ���1�I��!������)�忸e���1%M�ͫ��Y�M����������1�h�,���&h�����n!ebBweI����cF�dc�]��^k�x1���+I�F@ȓ]ߠ�,�*
����t��2^K�lPv����{R��a�K�� �T�R��&d�O�{噽��K�g����v�Byv�I��/)/���V�٥�nX
����������cY�`h�r�n-�\�WG�A�.:����� |]B�
�g�N��?�T;tHf��gM{b�}�hzir�����]>=b;v�8d%��r;O<�e��#�z�l��!q�v���N�S�Hq:��rp����<�����f:%�}���F��0myN��\H<%`䮹����,�~}ST��g�uu���Ϻ����,'s\����"_$1>����h��>ڻ��Ł�����I�"�Z��}>=򳳳qTf�al�O��K����
�qp��'�Ѳs��$TaZLe�Ҩ��)��Is+�يx:�Ǘ�{�Ոx�-�bk��{*2����&��4�dHb0���r��=�`(���D��ӧ���W��kݦ,���}"4WEi�%>Sy��u�e=���u��}i޻o_��2^fҬca�-w��}_�~F��<�g������gΜ������C�^�6)5�:	�K,I�H\?��������vN	B��e/�'�u~��dQ�}j�j�J����*���ڼ_.k��꾵��+m�-L������<v�`Ne�9;J)N���F/g�oP�ٰ�ߖ	��t�Ѩ�)�t@A�2�P)�0����ô�u[�A���K�?�m*�#�@�M�Ux��ͼU��;q����1�\[��B�@��Y��o\��H�؎���0��#Ii�K�g"G'�{��U=�h�Cv���PM7x�6u5.���ܹ
��,�� �\������4sብK.Y�Xx���%J����ĕĩy3����S�o�{1�c�u|�q/�<l���8���1Ӝ��c�#^=z��'�R��1i�e��<�]�%�9�"!t����Mp|g�6syL�e�\g�s���2iv3�JU�$�(��^7�:�����t:u�l6�Nh�z�<�$>��'�ϑ�*���u��ŋ�.�!1bj:�����r��;$$r�x�O��3�؏��c��|�)�������L1+��%�}���\�����1>�D��t����US�s�7�y�����*K}O�[�Y>* Aa6��4蚘������G�9So�`	�3�ʸUL���a��bN��ρcI��C�_ZO]]�m�c��m�mف`y/����s���q�#���y�����H#{H�}.ٕ�_�.� �����h�D �l1]�8''�F����n2r���Lz�A�������2��#��L�M�����;&!h�����$��$%##��o޼�B���%�_�h�c����2��O��>C/O��"[�I�� �@W���w��k��RJ�>S��K6���b����H��!6�=�>���������<��N�7D���LI���L�Q��?��",VRNXl>3��˅�esC���^k��p�MlX��h�D����
�Dl8Iג�𛾴{�d
*KM�*5؝XAA�UbU�u�R'�x�pa=�	*�zu:d$ɜB�KIM]sc�#��i����7"2����F�R���)z�y`;��K�w�
O\�<����Nu��""l�>�+qO�����Iԧn����0�|!'����
*�T�C-<���a��yDbLA(��j�c�J� 2�ܟ��ݟdbB�0��|����48���w�;l]�e��%/��������#�����?�q�R��g�-C��H�m��V= �������PmO����=Ω�����	}�ɐ{�&�%�qa����赹�P�!�R���˼G�{N
;/��<��Ď��am�a��]J�2�(��e��aB��^y�]ys�������h�KPQoG�X�K���]���1a/~��b5�� ��Z>����'� 0|q�S��ۉm(y�FM���8�������pI�mh�ak8_���$%-��f�\^�����o�UJ+*��H#�=�W�Nj���cr��$F���BE��$���܀�5���;��4H���'NOB	`NȂ���ƿ\�������XȌ��+��e�v�֧Gě�kC�L�z����`0J333���dr�m$I$�����ǚ�މ��p���W���� �ڊ�����g�ӓ�����R1��� c"���k}I#�uC3Ő��b@uf�ͻ�>;77���E��x�s��Z���Pc&k
�{H&�Я�nddęL��C�M�7.}�I��K�DTh^�,Uc��<��LK.U\�������,p��]�['o_z
oW�,[�5���~Jd��x���Q�m��<WK������&	�O�BY���ӳ����"¦W�䭴!���G&I�ۻ�����#��}����	�_;���bZ��bI�ʒ[DG�t{|z��qx���� f93�J[�P-�oK�i�{��俠ĹQ��w�`yaA�d_� �N)SVS+~K�඾�;hyR�*�U�M��d�#L��'��?� ��ԁdw7DU.��f2h60�nY�u��ݎ�jS��CU,�?2ݵXW]7N��~�5Ч]br�n~%a�{������PW��c'��KߒIJP�B�e�]8��XM����3�溱��lK�m�_�
Wۆ���M�� +B<�<a!~[��\02˧' �l�V/��nݺE#XgY󔽉��U�Sn��~m�nX2j�1>f�Bm���)"i]bv���%��֪:%ޟC�Ҕ[�[�[[�#JP���sRo�AE���{�B����G�/�fՉX�%V��fQi�B�U���0B1хqH��Q����b0����ej���- 12�I���jH�x���bJ`��nc���{~@�1��T�h�@��J�Zh�)jY�s(�Y͓��w���;jp��-�
Qtv�G[D[`%�7y�k�vuu�v�e2��ϑHM��d���qq����	LH5������.�q��"�~#n�@����'��}v������;d���P�X(.n�P)�}�E��TВ+�o�QUU^YS\���Gh��UN<x��x�[�������!��t�b��~�[I�����8`S�BLu�Dk�����BC��j�na�}�7�T��f����0$�Q�'���ږm�����!}�|HȪ&8��&���	.|���7u��3��1K���ŚJ�̯5B/��x��B��(�98�������1��R)P��c킔��ebl������Kv���B=쪟tu��@_pd58[�j[[ۚa6 ��d�Sb�é���
~��f�8%;����g|���ʙ����ՑU��	|E��snDTTU�ޞ�[���ñ�����RSSS��Sgb�����6�����4°���4$�pWG�	�./����T(���S��م:qI?!��'	���gϖy�C�����!9�V�I%�rg�!Y��:��^������`0�+���%w*�~�
�(Om$)\��^���q��@Pb	[z�]�Wo�o�u��Ԟ�4�NY��\}MESs��N/�C��
�V�eH��ܒYi'�(R<�l����N���I�;��}�a���;`�pb1��x1��qw�J�;Z��-48\�s1��~��?'6ӹ�Z查U1�U�'$��F�0L�����i���"�Ɗm�s�1���پ�n�p�C�/0��la�YR��I��^^�MR�J�xd�)�h�:Š��$�N�n�{��Io�RS���K'	�HYz��b���Vm��z�8�t|�d���\M�ޏ�׌�>�mM��s"� �ݤYy�|���*5od���]����I��v�Cm�1w	������imm�_�V^�cf=��W���g�b�Cs�K�)ZH���������Kh�}H�*�˛f��-������_�s����B��d� �<F9O	E'o���5Մj	4�	t�g��C�,�Ǉ������{�s��GbccG��ӫ$�g����^i�Pȡ��QP� r[ab8ͅ��v��%�.��	�	�8�A��$�� .�0;�	C���Y�[�_(uX�""�pN]m�'r�nc�MP�uזk�N��u9��j�y+�%;�,b�q��N�,�`��z����2a���$�=JEX��Wyt�Be��P3�e�&��÷۱��dKD��m��F(k������4�1�L�W4bQJ8d�v)ʥC��\�n�~jdj�P,��j�J"�^XeC-�H2�J�_��]���)Y���)U~l5oN��%x/0�X���@�Ν;v�Z�.�Udv�xJ�bmmmj����R'�W|��nag��&��-j���+�%s 2k��);�
v��?w�������~F����!�8jU"u� ��������{u{��gQ�G��L�MY\��Yh��Y(=�����z���g���G���7��$����%��y@�T��h�u��^�r8*�p�+G���*55A�?�)'-�Y�8�=�R�a�2IMZ���>��k����^��ӓ糭&���W�9��kam]х��$��ĠV�h���\�FaQ�����ur�X��1�CR��������I*6%�Y�=;�K �K��~������Eз49B��V����Ntr�x}�ZY>��/
s�eK�"yv#Iv����D�#:�ؙ# ��2�;�	�޼	�����X����b(Ƭ�\X���x�լ�hr�9�7oV*EH&<����ޞq)�:��>C��-i�FFF
���
��#��\��Q�����v��	�G­�j%��oxe0�0MMM���e/�+5�^�������v�e21���C� �,����nk��������]o݇N...1>6��~"H/5�[�cBFmג,�y�Z2}��x�sss�fD��H#S���T���������)��7�e��gI�^�F���)		��T��ߋ�X�C3hî�ҶQ-+��:_v@M�������atnoI}��J{�[9���2��(��룃���R/��*����[�(��#�����9ZƤ`lR�(�l"�,mw�X ��!��ۯ$Ƌp1]m�}nt�6V���([���$\q�]����ƈJ�O��3N�#��S��r�E,t�E����r�%���~gt����#�:�ʆ����+�eQ����
;�a��H�Z,�%;�j,�k� �����:H0�rEu��ƶ�d���+7��f�/�|������<�����b*�in^��*N�J�'QK��?��6]UzkI[lS� ��9�|H����h�9-�;Y�p��Z2�E��\�-�oj�Ֆa�[���DH�^\S�T9������߾}�"[�k���
q=�������~m	D��T�v�j��7	�.d�%P�@&;Y��9�dQ��4���I1�D�Rv!�ц�
���e��U[���Z��AQ{�-����!9�Kʒ˿d�`���,	��Ҝ+��%8���<�V���͒sx[�y?���_I+Ÿ����-n���l=@�sPSx��VBBBs%݊�v��� @��/��3l�4�FGG�b�s�(oǠ�����;.���$*���Oe�K�ٚ�Y����E��:;B��I����Ҋ�����&�P��B*?�9���\�ijrJJH�O�h+T������䖝�~VnO��CY��=50��!J��]������>ZZ�T���_�1�(�եEa�Ɏ_���H߃�X�Ш���0;���t^Z�Կ]�݌����N`�H
�tJ�O�1��-�΍ַ����TX���:3��+	yj�8��T֙3g��髦�o�Qd��R�F�gI��[�1�e���k��*~nRtb'��l�<��P�-6mK,����[�����+�4�dn�m�La�a-�SǫɹM9!X�I"���l.��R�����R����X����KLL��~E�֜�pӒ�>$-j>�.-�)n��(Qg��
ǹwj�����i0ߚ�~�i!�������T��q>Ѕ@hI.)��������� W�5��mC��!�M���19�M��N=�����ļ��WYYyXZT-��ʮ�n ���\�	J�i�a�8��l�Tm�r���$�����������#��-�֪�¾�f�l^mħ;X{��1�E��.{e��.+i~��*�zA��"�;ˍ�pPZTBe����ˠ?���3ɩ ����Ą�%\�֤�y0tY�1��cWV��'��<Im�4����:i@�C�f���A���a΄{"R����b��,����ו�ħ`mF��o������Es�X��Xfd�q~��+>%D���f�@��*�T8�.����4>�/ضm8~�U�S�!�]Ju.E1'c��Z�Z\|�����!��F&�
���TD<8~z���������)�m �����D��o���_�����me��|��ݞ�[$'�c��ܤ�&����`��1�]��ɈW\�Vx#�7���<Ls1���$K<{��s�ja֓��rqq���X�\�5�Kb�.�^��#/�/��K�8F�^s�>�i��O�4֩�ޚ\����i��*v]�ܝ��HR�Q��k]^^��<L��}���qP=�V�~�E�d�+�%�P�=�0֔�)d���b���t<���- [dEv_c`WH����(�t� �\X}��_�E�q�N��4���w�SL����33~�J][)��NE���lX����֧���ws����șM=�m�,�Z~6>>�0籌B�n�%K�9(aJ��+: �uO���}�.v��c����gϞ�D��܇y�s��RYի�&:��)Gͦ!�W����ڡC�)�ű�T��T�mT*՝��,��h�700��Q]�eFa��|V`e/�ZcQO���,5�rN�O����ڞ�D$��WVj���V�i{�$��*���V���2j�I��[�g�-zh$aj�q����q<�'��a���
�Q��e%6�<���Ȗ���ac�vP�40,�Bc����gmlV(<
чp6�����!/}�$93�<�����\�df)+X��m�d��z����n{�m0|.a��
����	�m�g�v�|�tg�u� �@���T�-�@V*u4w��΃M�41垬� �kӚ��]M�5-�҈5��$E���[NU{Ѷ�����!!�w����A��]���W�r��Bm�'�3f_/MU�y��Al�����z�sÛ��mE'n�{RR2_�Uom��KIZ��wh�k�!XNpC�e
ym�M�jh"v���EEs7�rt�;&�u����q�t�˯�h��⯬��:�61�!�u�0�ecQ�RDć
B�	i�����xGNW�����'�פ� �hZK�aZ��H�ކ�ZV�b���H%{7���O�qR����n*%�ڧ�(��k(S��<��:�1����b�9���a����D�P��7m��^�c[����[.|����������;�tO��}R���W��}4ͥ�1�y��6�e1�攕Y�v!#�vF>T�� �Э��Èև�{z�L��(����X�a��U[o7h��hT��9'6.n�j�B�����q�?8;F��}E�r8vm��v)�WǶ9J�������1"���kn�w�{N ���;����U�}�����*)����&�<��� ������mܵ���\<7�N�q��.\T�8C0�疭�H]��a���[XZ��D��ș��.,���3��U�!y�b,�� ,Z��@�;"RM��r���t��XFV�8���F��QJ��CK�ߤ���W�6�
]��&Da�	��)��
�Rh���`�u=wn��dc�e�ht���-�Pgw�)��*=�T��z���>�&�
�|��H�����A�O��]WBւ��Bh��21��}}k�m_�Uj~���!��ݻ}���į���.TS���d�|�/��n�)�T_t�̼��e��Z�&���� ��{e��>��W8��y�?:pq,C�֭[�
7۱yd����ҽ�|����n�i��P}T��0��ȹ�����<vi#aii�ҧ�tO���Z�@��������6�/�����I�
r�����|�{E�k+�TN���pyW��:3�rĭx���zy��	T�? ����L{��܅��s���#�Sx2���w?|�����!����bA�\.7f���3z��ҨOy���/�|�Cd XH	�rd�߻��o}n�Dh�B#f;���<�m�>v�+���1?�,�MO��ϘB����C�Â����B��@�쬬�r�GqAZ[P���5��^WW�w�T��g�����iYY/ٻ��^JB���n.r�rV?ڐ_q&v�=��ck��+q���8��!�ؑ��� e4�G �Hvҷ\V#��Ei�<�;^sS����0���E�*�9���"t�6�kwC�7�Pa*a��ɾ ��J�Ϳ �5sP���K�&����Z��_��T��x<]�Ffw���SPV�h�d��y�L��iTT�!]'��EE!D� �=|M�^�F�3�3Z2v�����E�.���k9�xc�E�6���@㇕��ǀ��رcGo�7s�f�7?"�t�^��2���Y��A����%��qZ�*oS�#��o=�İ�!�6�����5��÷>� |�CIpD��34���#�㦩Yv+��k�-�P6+)ˑ@Y�.�"t��k�YY!ܷ����yg1��_Q�����do���c��k@�r�����#��*�g�x����(��!��X ��I@v1T1��?�v�|Q�`
�,#�7��s�ң�Nw��`~��鉶�����&�V�D�Ξ��q$1���tQ��bs�2̞�#��8�Q�M����}s��7C?~�,�ɇ�v���{�$"e�I|l(A/�+H�5�0���H%*�����i�"Tpk�YпԓR�������y�*�qm�wC����V�/�~Wߔ�^�Dχl������+k��h�H3њ�=�Ն���;�m;�8��"vJIk�'B5O��>��r�F�����roo/+1��>vUVV�C��y(t1Ȕ�ТTb)?�X�>��/�1R���M����C�A��~�IU��N)U?��IU��0E��w�0-~�I;�G��Ht�����D	�ZM�X'UՂ|�@)ׯ_��\4���[c#���w��8zp�(�=�@���߭:��6bO���� ~L N�$x��o��u5��Xq��"�f�i�q�<ޕ>
���y)a�.��K��"(����܏+��uKE��nbj*�K�P�⵿�^Yٽ��j��R?
BaJ�根)y��n�m�		��;ru~��ч� q�d;�7�+p^sƞ
�����ɟhҪS�<��3Pc]�]��"H���,�����y�]l�0I]Mc�&�������2�6�5U%$$lC-Cg�h�>h�M]�r���]��"��W2��*�'��{����k��S�f��>������#����q����%��&P������v��j�q�m8���t��A6�1	�ȣ$0�k� � uL�QKR4�OZ4<�����O���)An)��Wq!�璣�P�J]��%�v�g��~f��@'�Ҏm֚���]�Z��%$�3:}roȗAm���oP�L�H~S��*��ATUBowHMM�=A!��
�sI��&6=tש�v��}g����՘�w�^�g
Y7���ɢ*����Sw�c_JA!����!RJ��5��prhp_�����Ss�;T�ަ|a�c��P�ڇ���8Ek!g�s=���n�X��\Yi�� aC��+��K��3vX�x�����@b %�C㇟p(�9��v�5�0��i	Is�c�5(ot<��f6a֪ǧ5t,{PalL�&�c	RTHu��k%M�6�&&�To�,��W��v�[*&�hy�)��C������)���>6		��h���C�)��� �AB?g�J��[�#G�����Կ�&s�$M�Ѣs@�U�]���g�ቶ�J<^H!	�ͻ��Z�!/g`_I�����[`��y�&7�n<��)z��e=���5szgL}3$���-��׷�X����	�u@�'n);LL
]�\Nm��4�y�N�D�"Ӏq���5x\tZ��V��@u�N�"���o�w�����]4�K�_�C�n�~�$��C��G��w�{0M聺��N�V�>�
FH]�����G��U��@L�A�22��*�e��a߼y��ٳ~O�X�S�^#�TTI;�k�!��@�¬,�7�q�Q����.AR���Q�75��--�2}h�3�Ɏj��prC����N��	;���^j5������j=8�Ϛ�+���`�PȊ�?EG2x{;�9J��+9i;(���7D?*�1QRP�Ґ�"�C�5�k�C�r�K����u�OB�)�N�������3I��Ê�X�W�oA��j��*5�a�����D&9��g@M�����V�1>��¿�zHu�,/��/y�u	e�I0fL����M5�˗�����=��_�e([YY�^Nݳޠ
e`
���Ƽ@�f�����W�˚�N�A!��j#P[ͧ��������`	�8@�8���|f?=O�ޕ!������&1=Oe�?�YsI��%����C3�_򔯌��T�,
�k/b����Rg�v��r�Ip�;x��*�pr;��\����I�M ��GyB!y�s&y�U����V�%?U�I��;��3�E<	�nnUL<�&�:�R�0ٜ.28p�E\�/;Hs70�pfF
�G���/���=��ZM����J�M���};%���\�s�v���\y�������;(c���7�w���*$��>�����֢�[0�=S���8�����2�TtJJK���=�i�W��W���F����!)����%��峸�O��L��MLZM�N��(�_7|O�F�n.6+�W���4�L&�I���N��͢X����"�,ɪy�{J�E��Qlc�R����d1ؾ-� !�c�@mZBI�\�m�f���7�G��Nه�Y5��@�!L�{r�K%��ǮVi���- j�	���%�Q�
A��D��ֈ�
;��%1T�tM*m78���(��߻ F�3~At͍%_:Y�4�������^pi`I�JU��Ϻ$��_(i<t��6�哑-���a>h�zI�M�87+k|ѽ���'�<�/�+I��'3�M�p8�I�ڑ/P# }�����)�(��(D;jkP��pc۾ޟTU�7�UZ^�%��0��}�3|=\��`��i�9�Zt|��-쁈̬K��7h[ ���
jN��&��)٭�$�~�F0�'���5��}ȐI�f/P�V���q��D�� �<g����)�,_������w�
�9H����E�?!4DgI�Ez&�4��,��l��ٲIBo��/=_A���s�:�wcT�)f����o�E����Z�:���;h���D�����KlYN 8b�qR����WHc�����J��98Db#�V�}q�F����w�%�K���<j+=K� �<�k��f����(���h�{�#�VU]	Y�Bұ"++���q��d_~U�ڵt α�c�SmЧ��| ��e���9��P��Z��W�2=���*��DaE;���$�����h���H����j%��~6&|y�]�܁ۚF�[�$�lCW����*��&�-�\���K�,W�	Έ�ה�� �ݲ�?�&����ҴKQ����G�+��{���#��XuL�N�z֖V��xIk�p8���;�G�� �B��5��N-��J�6>6Jü+i���S�yh#h����l!
+>��(Ƞ�z���(l�bfFss����_�w�ٙC�`!p�&X
��ZsS�����աV�F�)���茏��)�K�8i���[b�T1�\��vY%�tS�MW7�Z3Y���t�:�φ��Aho����UMi��k�؀�~��������
֭��]G�R�A�p��V�N�S�?�����e��\ mŻ�}u%��]�͐��KAy
촘���X�������R)�h�����Wz �z�6�G$B��ԐFe?�S���</�UrR�$�C��kL�o�%N]ۺ	A�q�?��?/tuy��vH������t8����=�k%����]]ށ����xf�yt�d������'}M���P��'�:kɬ�@iʚ:-!T��)�`)d�Ql�k�H�̋�+��N�g������	V���3�	%l�=���99�W�>73��#���:;�|�9���|a�P�T��)��)HD��:��0GƹMI$A���5*�v�8�<RWW'lJv��i�íz-\>S���#����^~}���2����?�9���Y9�����O]�8{�s��=���Ͼ���F_��"���-��P��ySS�M����b�w�=�(ľ��� MX����Ɗ��1�a4���G�L��*�q<Nqś<�`x���~�ώܺuk*��XU�\P6;;�{
�**Ts��`���=׷�O�w����ѷ?��&�/�.C�[5�����ZY���z����B��J۩ۃ2�ON�*���Uz������Ûw_������!?�u��6�:���7c��"�s?���+onk��{܁���ʏ� ?^S.a�V�p��8ӕ��`�?�*G#���I�Ckk��x�-am��QT{� ���;a���+�'ږ+%�D���q�c���G��Ro�/MOLL\*�wOݦ\2%w�����@�V��B$��X�J�S�������N{����/�|0�x^�մvC�c�;dVxٓ�m��T�oKB5�yb��
m���PWE�?���������U�G���R��G��08���<��Y� 1�SPP�dZ���V��l����z"�&(�P��:x���prr������Mrn�������(=&@&��:*kB�'�ee@��l���e^��w���ڲ)&�i,RX��i��d`f��Y0H=�oG�y��Գvv��< ��}0�c��`��#�SF�~_�J�L9�^8VV�"��@�柠6ɉ�-�E=�1�
��O ����R�7��Z�=���H�������>�bWW�΃'f�$����'�̴�j��uh��]}}k]��GT]o%r?>!A�ݤos�O��k'G�>I7�.R�����<����d�v�i��.��cj6��$�gɤ&e�/���o�x905�F���.//���:j��8S��[{���R��@R����b���U�;]Gܮ\ܮw�H���ǋ�H�޼��t#]�7�Y��.BG�Ð�Н�񄄄�N|���\�n��&c������m.�
^�07k����<��|���-��[*�#׆|i`��
����q������4�9���n������埽��T�
�r�5eؒ�^_��P�kw4b��o!��ÖtA����J?�v����Qv������+q�LR*n#�wc���R?�@�T`�Wg�������	oF�PN��l�?R�p��xY՚H�=Q����၁�&�	n��}׵�E�FMTs.t�=��C���ev�B�����.�00��;���' ��KNN΅�I���f~@�*l�Z�:�-u��T�q
=@�lto���:5���;&�0m�l'@�	�md``��� �����������SS����k��j��N�Nnb	�ae��E��a�L&��E��g��1>~LPu)V8�(���i`�9��e~~�1r2��2���R�2ۆ/���m���������Y 6�q�2���������h�()(�}Y�j�J�;-�C������p��~�e�*풖^�#9�-m��κ�|[	������:j�{zV�f�*�K?c�*�P�
��D���N���x��N�f�هYY�ֶ��wp�S7s�oٹ�S����7�`�[3�d��"���˥ۗ���6v3�a]�ͥ尸�J7��_T!p���Wx�S���/���߃��A� ߴ�~�~���Ļ�ꎢ�R��J֤/n.n�S�5>��x������)���%6N�T�5��׷>������[���v�Z����~:43_,���7���\�gc{���\���l�zc޼yc��x�L�`ȅFH!b��A&�z��-���:<I��O( i�f�&�ʮ�+�������8�7^@E�3j]:F��,)�\�w/++����L
��g�RySSv��Gp{)��>�M�n���ra����g�Th��z�����p�2��'vs��Q���( ��]
�4��@�K`T&��,=�/,�q�̬=!9Y�o�[f��^!�Z�!��D�P��"�9�e@0ʨ#��8;[�����q�.Ģ�x���r��ZIC�w(�`T\Tp L@�_�e�;������,��RS�A=%x4��6�� ��UGG��7z��Ϋ!7����(r�^��Η���従$j���@5a�s���89��%�VE���u]vϵ�v���o���������m*|�|��@
%�\��ɹ�s����֖�I��#���ۏ�
E�2�( Mo�;����{�֢ٓI��ɹ��	ߴ�]HLc��kT#H��_��X,j����pQ=�h�:^j}s�c>�����%q�e<P��!�Nm7C�*���7�M��ǎ���-�F���Hz����O�|X��i����?�]X��%Ĉ/!�B�{��D��f�Ft�G]Zt-����o��)4�(()A�|��Ԝ&���*U`r�]'����Ꜷ�y�F��/����(L�gtT���\��o�yxU3~A�Bc�����	����^��Ǘ���=��*�i���7o�PB�k��zY������5%�O���UmcZ��ޏ�9���8cTe�+�~m0#��ѣ%X��N�a+++wu��K�����)A�\@e���nZ�g���B)5��f��[6�9f+4*�$E,������V�����6�h�]��\2��G
�e7� ��}���\ݓ�_����=�b�*A�u�\�Ţ�����k��İc'c�����d�y�^���#=K�˗�����de�z��/�qP--�ǿd�k���?����f�Y ;�o]�n� ^C�S�.�3�����s����z��]�N��qMt`��� 1x����7TRz>a���ru_�⎛O!�\o�����B����h΃D/w�o��l����`*x78�>�"6���f�(���/�.�^[rfHӳ�3#	��
�X�B�hgX>��*SXz�|x	d�q��ͭzj41���B��zIS �A'�"ץ�M�%&�T���1�d��(v(�#���>�*��E+�r[�REH�q*wʅK��bb�n��*����c��:ǼW{�{z���jf컗�o��grK�8�# �ͺl퀡���_�I|"���̬	U�Ƭ��H�r톲r"(]��[qC\�&���_ x�s��t���h�Bd��P��8'�Nz�P�=��|U�B��om��U����^xx|W+:1U6��-�S>ഏ��>�A���N0�mT�K_���f�[mM�~ff�J�J~������*҄�j��P���ļ�����I"j=�HK[7��d���C}-��_��!ȮBR� ���1�� X��^���� `a �o��P�����FC�a�vY�T# �h�Glնa�'w����^"�Qӂ�tё08��×M�3G!aGBJ�Ȏ��ǔTz����GxrK<�Njj�������ȹ��?�V�ppq��㩂�Dw�+�>���'O�m�Y"���҅��C.�8��ff�P��PUUUj�y�,�Ȯ��s�*rE�d���7��������R��Ӳ����e��^�S㜛S�M���������5ϟ��L:�4o�1��&ж�(�鍉�8	���� ���ҽ�!?`�~�ay||ܝ�Z����r�G�e���vF����w�������_��p��Ѫ�,�}���v��[���ŋ���}�Q�
7D�?X�cf�X��K��J	m?
	}[���n=��u_�+��;���6�@Iǅ������-��x������@� ��9�Bd�r:��]�t\���u�e3�5���������7�ͺ�,~0 U$���TH� �{.�����;t�R�Yx��Eitr�����ߡ|������5�l��CzCV���h�;r�w_d�T\��Dڶ��ۨ@��Iuu�X]�Ԛ+�S�Uh�<��G�>�g�V��!҉<6��n|��h�Ľ��
Zp��n����}\ZQ�w*�P7�����\+���$a��,�s6�Kyk�q��
@�������_V������ˌ$�R ��)���kHj�$�+���q�d���پMW�9"���	ʟ���ǵ���E���J� q�+�~�X*�<B��s���^�M��gi��j 9�������҈*��oD!jxLd7�h�}8�|ޞd�G�(yo��9�l�ٸ$ݫ|���!1Й��I_	`�ūX�"�T�hZ�]t�fx��#�K�������`��U*�ME��>,R���aP�Q� s�Z�Al�P!H#5����j�*��!�"F�L"2÷�	������[�������޿��sεo���,w?H9/^�a8��x�fm��}�.��J��ߧ�5�d�ڷUy�Ⱥ�0�ځ��.v򣣣�٢`cĈ��]����{��N�/˃���+����N]�w�;�
e2�۱]II)B�v"�d���Wɴ���E�y��JX�x~�2��n40$�J?Ȣ��&>W�xl6���,K������_�$&%��W�4������8{�t���@���ym۽���/?)
��럵��T�_�<�d2�@�ħ�*M,��h�q�̈'�>ߒ�-�p�&lK��폸�I !���2/�u���V��S�����_�ۮ�V\R2o�TpP\^�����A�?�ltp�־���zW]&�@rE������D<��8��6-�%O ��0����[����By��@�<��s� �Ո�L)�Π�����|ЙA��	y���`�Y�-�_�<��7>��x��7�h<X>��I��e�2*�v��V��Jv>:�序P|��ˣ�.����M
�\&�UB'U~��oT�/[�tϓ.�C����|��T��`�����y{���B��h�'�N��\�f��ۢ)���]4F���]�qv�;�Ν1؛ׯT�0<��K�7���R8y�+$�uO�����腚���jY��@��]A5g��@�UcZ=�ؙjd��hxm�� ��W?R���I�0�S�5���F~�}�*_Yf��L���W�����>�F������+V�)�%��Krf��.~���#y}��N�:�E�K�X!�o��Hkܼ�z�Fғ��߄�9���>��zwlӹ/lW l�N�a0<�xh�f5�}L1;xkY��<NFG�t�Z����s��}���w��M�0�f�ɜ�0�8O.Ȼ�y���������ߘ�xϺ��孻FFF����|�2�`�)�`��[�PϜǕ�9�Kw�Mb=�GQ�G�1���*�TN��I�rURa�щ�gt���ڪؑ�)xz����[YU5¤�]��O��W>Ag�I��~�.�����2A�I����<00 (d�k�dP �9�*N�:���$`�C�Z%o Amu4k�VU����ŀ�3ʽ�_k�<��bY��GGL�g�]���Vw**f���X�Ó�'>��֦����7@0�D)��>���ZXX�j�ÆWY�]h�x5�>=;���AǺ+;cG>5���E\��a���w�Qr�p��\�s�u��ѵ�ׇ��U!��c�Ox� -;��6�~��;��+���o޼�?>>>�����rӉ6&�\�J�p�8�;-�Ǎ��/�1`�@�x��&�_]�w�ch�����(�oQSS�z?����c�[o�2ue�� �z � 4*�Z���t?�|�qoPಟ �[��IXw��;��܃�S�����ܪ3T��7N��i��k�6e�U���H�5��� {(��\>��bW�.��hO�U:+8��\2���9�n�PWIee�Y�Թ�Nw^�����@X��lu���t�p#�!�2�����(��ȿk�J�����9�$)�[����p/I��c��ٹB��H������79��x��&$��Y����]�qv�xOϰM$�GK�����o�r��n��R˄/�T�u�(���Rxl��]P�dY�z4�MHѮ�4y��	��+5�e9U��:���{Co���$����B�C6�%<��s�஧���˧zF&���$(lɘ�ק@_2���#�;�-qT�F<�+u��5c���!,�W\�~���I�:m' �/{��$f���F`�@���O��mc�����)3!n�:[0w=C~3�j����Y]Z��3�
z��ձ�����.<�������w@���-Yz�{��`�kcB	�� �T�Hk��Z������2�������O"��C@k���ܔ���sލȧ��0f���y��j��T�����5�k�u,�1}�SQ��f1D$uǾ�� Cm_����HNNNy7�J��D�%ݥ�?{���
��� ���Ay]�^����3���r�P��V);w4��ݒ��.��p�Pk{�UYVZzV�݃,o4�=�j XiL��H�m�B��׺�~}�FkFo��Z�Ж�	�?�S�5���'���wSw��ͭtX�9%��l\�ٛ��"+g6�O����2Q��
�~*\a�I'�5"�d������O��U�����)`l�/�+��8ŞT���Z�́	�?N���A�~�R��
Pvっ����q��y�}�?�R"GEA8��C�C-q����.������ʈ,|�NO%xɻ��p5�k�Ÿ]��+���Ԛ
��q�#Ną��8��J��p�N��^�y+2픡�Ri��S�CxO���c $
ۘ�i�7�Y;q\���yFS3�WE�.pK&/���:��^�,�\��lܮs?fu��� �Ԉ�\&�B1��^��a�0^:���;;�8Ac���0U�z�j	`,�m'�W0u&0� W6X�
b�K�������
��'�$�nm`I����W��U�P ��˄��0],	��K����ޥYd:�5
S�^+�W��H���]<��:���S��x��F�����r�Z��p.�Ķ� ��ȈQ�צ��n����B�{�6�����X�@�3 yR���Kf��XIWxCW��" ��NHagO���P�E\n20�%.w��Q �=ť�� ֑iހ�22�j�A��(�K4��^O)��w8��][Z�w��5K�������^�+Q9y�'���������!d4k�j>b�!688���N��;��.ƣ��ʀ��]�z�,ʉ'�v��7Y}tg��~�3k43�q��F1�m��<�D�R�&_ʊ�Z؎/�X@��܌�|�;�`�U�N~#̮D6l�y_����
: x��g����E�k�/��ѫ� �i#IJ�g�t���Q-�|4����ҝݴŬ��,��lL!lT'�;:f� ��A%�6&�G-/��];�G �l��LCD
		麨����S�W����8�pX^��/��H�Ed��{�A��������k;��	�Jգ��Kh����Z�3j�
)�@����a)�(�\0��\�氞m�S�6�3���q�r�A*����.�r�q��D�&�� ҄�i2���O�,/lo9(o���<���+�#�D�� p��<`�+w�}r5�eq�S:�<�*��l|� ��o���Q<d��T������������{���"<�j�/o6RĲ$�V�i������V��h���`��9i�	�fKQ���Ƨ��2���077'��[�w��;�K�hV��

�����`��q�5}�y�v&�LfB�>����{Y��mɺC�b��2�����m@�E�{��u|�/c��4@�ં�'3-Y6�5��*(�8 W3 -O\��Z���	4]<;z��g��BI|�m�B ��r�3�o+���Hmm� �fڟ��5N#p󼩗J
��	
�1����|��?�����v8�P��*��{[�@(��8T����A|�M�������@	/"�ޘ{�BK��2}%1%���?��Ɍߕ!����F���y9>�
ɓ$������-,�� ��N�-����K�Z�!�p4�OEiH?{hq���
s�3X��Z�F�9�6;;� U��9~؂�a�3J��o�*��ۺ��b����0M�z�e��5P�m�I�œ,(�Ҳ�(�m�g�z�j��!�bV.`0<��rI�)���\T8)��
R�Ѹ;%���x3 g�x�r_��o埫�Í94�Q*���:�4�*���p�zO�);�zf�s�<�d���8�s���pxA�Oim���徂!��f�d3���Q	�?�w�f����Ə(� �/j��ʠc�!����K�/��3��^����s&����{+Wd ��̌��r&��gg�=����Mۇ�5�������@bo�ڷhhi+�.�(W�n�8w���� ��}f6�P����v�o��i	0����	��h��>�w��QJC�Q�- S�L}F�ȨQ�4N�gQA'W����|��ԽU�DeI�N�1������0DC�^0r�������I������g�52Q�mdʰ:�g� {mp�̒l�rS�m��e0��ٷ����l�j����7��w�ꉋ1HKXn��F&M�+�w��)�ş|���W}��ƺ���=�ɝ�T)��ow���X��|�s?/�A\�W5���� 1`���`�w�8t�a���RuO/?�u�4��׬���.Աpu���x���'ʐF3;lR���ɷ�~�m�����#���% l��7��:^wl߃��`dq�4��������r5�ߙ��F@��$�8����[%u� �O�M��r�U�#з�?7\�/�ٛ&Ä�B���J�8�lfY���١;8o�ܦP��?ّ X��fZ�2-�Z��C�S23h�����Zd�yǽbO!d�NZcԗut~�u�\��*v��f���,�ikM��JY�zi�U+p��O��1h�j�@����t� ��-"�=��8��e�����`�[�=
�%%&Wȍ��o)�`E������p�F�k�����������澒�bD�6]���4W��;*G�vBD�l,ٛe��/ٗ�����	Q��J��R�@�f劎@b5c���@7g ���U���uZ�2��2G��Z���ۋ�gkCr�&x�ůpD�S���*�eP�{�;�i�R��N�8����39�� 6w��T[�X�<���h@t�U�-D�6��ig����� cm��[��h%�Y�����PU`PЄ�e9(g�`ߥ��:(S�y��U�nԦ��]%��˛X�i�����սC�����:�U#�2�j����L=�oMߨ涁�!ո]Ȥ���	�P�W��+��o,7�ڐ�M����UtU��`��%n˸ZŔ�X����+%��Cr��@+�+.�'����ٙJ�G�����
=��uK^�f��]m�֝dXi��1���o�L�k��ɿ� �b�o�B�}T�}�:T͞7cmUW,�8P�e�� �5�kL���R=:]}�¯#S7���=��3��kS�l�y_ ��� � �RM�@��d��$@�VU��i��,Q���8cy�wo�$xI`�n��AFe���F�"������k�_�㌙�]i_s���V�;��B�}���O@���������f��{|���#�����K��@dzP�eP��A��WY�� ��5M��HW�뿧�D� S5.8�{�|�/,�Gv��FL������s�$��.��Oච��˨�im|L��O��6S9�elA"�]曃c�8����u��8[����X��k[�q�@@h�\&c�9��T�d�.��OJ�.�5(G����\��Ayǳ`rpa
X����񨑾�6�(�ց�4�䷟�Lf�o�Kt�M-U�9�?��ywЦJ��B�W���ȭ)��n,��o��;��a�jJ��������]e�J��N�?�a:������0Nõ[��iH'q�����R�%�2d�6����L&D��ލ�.�ut6q>^ؓ�EO"�#˛�V�e�����,��8��3��L��o�3�޽{�����͠�KQ�X�1�X�t�����?����S�G���T1�/e��u�-a(k�[5����nH&o�5kB7���L�,�ލ+�B�?:��zyz���&���b�>��>����
 Vv�r��*�����cu�rn6�7��R��N���������8���>+�)1^���3������R�,N��df���X�{�R��hз%8?��k�;qa&(O���@ؕɖ��p_�K���ˠ�e��'��!�.P� ���U_�-�����TdzB��.�I���d�ŀC�R���@x%���k���M����N89�U�iD��C�X�s۰��X"��@�pޠ�����v)dq}�~�X3Z4�f?����������EZ�W�[�ٷU���=(�{]��Ş
tn��101A:��t1ʍ��7.��):Gܱ��\�^d�	0S�=��^�&�9���[�Vp�\ɸ$�P�mg�p�^X�<ܣ+v H�J��rGg=�����Iw���2�z�����K���n���ۮ]�N�?_�]U��Ot�SY�]�d�C�������@�q���������Z6���<t�'�����T�8բN���,(U����O��@`r�Qx��<\(˕.���B�[nL�$�Ȉ,�MY�)_�mh�P���x@�8��dq)o�ӛx��4y?`|0��|�#�=Y\�~���ӛ��)�M��/풦1v�1�˕��t���]��1�䷒DD(Q9��U-�Z����r7��FU8�2bG�4]0���0�W�}��wO>A�gZ�P^�!�L��ч�3p���z��9vz�ja�Xb�,?PJ
+3um�F�bT�G��>�����%r��� �پ�Rqy�t�fm�ї��	���咹6��%`���1m;�-E�M�ݎ��<�h�x*�݄���b�J�H���3���=��%���zkd� �!�ʤv��=�q2�z_�%��UŌ�Jl��s�kI�tS���b|]<�M�~Z���k�!�ם?	:p����U8ܩ'W77�B�q봣Tq�eb<������,��T#�P�>�|��B�,y��%��?BD�A�׃�,:�W��-琐ܔ��iz��C����O���(���t Um�R C�S��	�3��,�_Z���t`�{���2�/^%!�2��U��j0��������,l��s�~j�R�qQQQ�(ϻ��w�C��s,Z��C�Cn�o�t6�	��K��`׊�����SG����}�s6�&hGr�� ]ɽ/�E�F��%0�� �D>���4#�E�;����8ם>Y2GF�b�����S�*,�w�u�mh�i�4"p�����@O�h���%���Ρ �1Z��[Y���Rh" A/iނ��X�0<��w+�2S���;�.?��wp�����-����@:�w>�����N�j��8�sN�g7��*���D�w�f�&3ە��ϖt�]"x�m����nC�}������l�|�WI9���,,��]�_;{��E���`��t���Q����P�<B"K===�k�́H!�/�(���.>Y}�Ӄgqu�N���:�e�y���7t �=��S/4
��ɏ��݆�W�ooJ�TV�� ���7H�q|���д�g;�`�A߆A��pBLg6��g�Yk E�@�SH6>��q��r6B�;��#(�{�\�KȚ��8=����A	��AH�@����qi��9u1�lrP��<AU���[�S �Mf�nk� ��Ni�~��K��?�߽y:a
]s��MV�d��$r�O'Iz��t���M�
�V���$J��lc�]<����5 ����?	϶ѥ���Ubo3.7~JzN\� d_�S5�b3N�/�� ��O��&|�Ɩ_<ZQQ�-�oA�g����᪢��|�FEH���R\��F�l��� �,G���p�# 7
������@���3�/q~�,�w����tj�q��_	�����괞�'B�7�9��Q �e�O��D;��\�1�	�T�C��r��m��E(9*U  �	>1�KF��d�@c���
�=faȷ�{f�]�0222.##s�&������$�IBI>*�R �U7YOrrrpi���� �q�;��B�9&�r~�LZ}��;#w�R]�w���u�L�?ԅs,�V���j������Y�^	J$�7+�	IF��=�ܝ��a��P�q6Ó?����J\��M�kp�%����ʸ����N�j&*���>�;/����a*�ol;?�a=�*�(��C%��o�wvιj֞�΀��	��=48vǖ���~T��Ķ�d����Z��>��Z��'?���/Nz�[�_6g��<+T%�s���h�p*��ȚX�sS��z��{�<���������w�w���ocj�J<�22:����︿�|~Dh�L��D��:Ď�Q���ju=�w- ��� :=H���c݇Ǧg��d֗�� ����:ئ.Z�CY ������9e��Ci���h��w=˓,_��7�{h�1�^7X�+R���-��?-a�6�TG?�Q:ՈɆ�������� ��d� фd��Չ�*w0�O�=�z�v�pt���gȯ�Km���U(;q2�����pk����W�;.h ��%����ꁣ�hu�����%�?�
���C3�DљNU�άt��-�e�gJ�2�?R�n�G������cg{�Z�bB@=�< h/��I���W��s�?�Ǘ�>�/���tu'Z���=YѺ�{5g'N|�q����8nI�d*eG���@�_�Qe���0O�����%@�p!�0厫j�2�!�v�w�_
��ne����fm3���fm����v�͘ni&#�,$M���m��I��)DK8��T�eԬ�
/�ؓ�a���De�8���u܍S�)���l u��y��N7ʒ��~JF	᭓d��Pۘ�96<�g����{i7D����x�2�D��j�S�rT1j��o�� �@�_,��i�i EdE?}��_-�ޠ�4)k=�)~�V��H���#��g�k�?	�1]|�U��~*��2k�~Q�M�]��г6���m�|���d(�,g��o���F�s=c㹣�ć|���͆����������o	-L�-��&�����ޝ�N�>�#�j���/i��u�����ݽ�\�;t���*��'�"IJ�����櫛m��b���?Nφ��%�*h1�U��b�����z���@͓֙{�:7W��w�E�H��O̗ũ�2�^e r5@���4|ZIy���|�rʕ�YLd���ލi_�;QmsJ?5����Î+�=��D�؎ѲkP���k�����3�i�.�ZE�(	ᓪ��!W�>y���{������ �>�	���H`g�S��ե(��sVo�ݾ�ŠJg�$@t<	S��vJ��G�Oij�/��Um�/ ���|1�U����u��g�S����o{7j<c�xͽ���e�L	��,D�.�D�y�p_����d��=Mޠ�೎��V�N��U�^4�P���rgձ���3Փ��^*-�*�!ֈg|}}9���N��s�G z���K���Āv�Ş�R~d�
����7s�C&dI�+�6B�� q�1�A�P�1P�}��V�]��b#]=��_ɳ���7LܱՁ&_�X�i��p� @����T���ů��Θ�<i7m��2-ŵ.��}�o)���������P�!�q'�3&��'��=(�/�RS��!Y���'MxJ3��}is�y�S
15&U�s��1��W������ų��^�-^'�s��~�0�Ŋ=���g��Ņ������x(Z�Oe��A1�{��eJ�h�;?�6.�'o$u=����!�?P���y�T�vtR6��oHk�yc�cPu����38sAO�=������-�}x�V'٬��ص�ؼ��-V��'0H5�Vi��咑�������y�u�6��\������Ş���'a|��58r~%��{���av�ǜ�)�.D�u�>ٜ�~ك>���F��L�5�6�������VVQ�$���V��sظ�����#�=�ʂu��gPpt)�-$uWR9��%%�ѯɔ`�]ŵ�^_з+����U0U��ԃ��[G�V:��׷Lp6Ğ��W������_z2+�,"ˌ�y�Z���U\@�| >�h2^��Y=���2g���;��k?�0���KU4��m�֝��]S	8��s|P2��;�!h���j�J:񋣠�*"��4�­x��g�X���ԩF Ow�s�2(�OQy��϶i5`�=����[��$&�Y�J��xo��ܐP�+5����/�7N�q�-m���
h�1�yC�B�| �b��kQ��+�r����ut���N5cH��+�g�ݻw����Z��a�	��ac�J�~�m�	t8y��3�(�����V;"o�fo;Y�L�`�J~;���[}�/_�\l���ř���À?~��Bօw�r��+���#K�,�W�ݻ0ݾ?(�]9����K�ζ��T�
, ��c��*��U��OS�+�FA�e�Vra���D��}��]1bV�x�`rj�T����L	���-��/?*���P.8�����u���Б�Y���ok1�'M�W�� 7�0
C�*(�8����7V��$�ʡJ�hr�X.����2}�eyy��G���r�e���1�6p~S}�@Oo�`	?��-9*��p}&�/c��N�@s���uO��X���4���1�s���}��$�(�/���2��Y���n*���{_P�_~��PP1�mf6B�y/�s�ؓ	�U�9~����'��ekJ�=����P�(�͏<e+y
8c+��R�nC������������L�_����|/��C�;��C�`�N
{���Ϻk�T4I��Rp��ڮL��X���"�Z�[Z[[M�P�$�,� �4������e�O	���)�V�C㝪�� ���wh��2��'ෆ;�,�Ğ|X���	�Ne��l?MN��~:`�R@s�բ��w}I�dsX����
��$����%C��JFMM-r��rS�'\o{F5H�Sr}S�k�����y�~W�ůs�� tl�>?w�
	���6(�~���Q^���!9�-r�W��3�޺����ҶJ+Fr-��%�����zÍ�D}��bG���Y��Ќ|b���MB@�#������o?V����nB�����,����ۗ�<�+ w�at[�Z���#	�����"���H�q�&S�m´
�B�{$�ᤷʚ53P�v��K�Ge�%AF�v�a[J�q�e?`����N����5��r��O��=���}Ͼu���H_|f�C/,�6<�\���F����Ľ�#�0��,d5(EhE
��7`�8 �5����I��m;��Rt�)�A�^�'�QL��%jTM�g�#�G���/� ��`& �(�U�ʔ�&T��q�.�����o0�^���_�l$��K��tHS~��zt�S��p�]".��	[�/��g���b~-cu(��=I[�>�.�v6Ny�f9�3(���`,�cR�ke/���������N��*���<D��>oL�X����*u�N~�	�cJ�� d��||���
#��iX`�sp��rT�$/��&��v��V�	�%�&Ը�~ɄD�%O8�_?�z�S!i��y�w���uLI�9N4.7E7mB�B�;_�t�9�V�eq��(�y�}C����9a���)\��l�#{�����+?�7�+��V��Y���-���y������x0�q|�vO�F˨j����;�(Ʋs�Z����w1��`1��[�b���Ѻ����LO�r|�����h3�P�ᜈ8�i�%��/qk���R�V5�I�b�+�2l:n�q�������NB1f�hY��.��/aϑ�W����tu�xP~m�̊��F�d��n�>\(�[ڮ&��ҷ?R�Vk�j(�2��6w��Wސh�/>a� �S����i<�ߟ|"�α��S����|n#<g��h� �:�:�yh�!f��z�-=C}��WP�����m��T�՟Q�-�;�僝~���>��Z����<Yh��T�]�������6��t����۬g+����o�p�XP>���Ѭ�@;<��zr�m.G=z^�K��ϙP;{����$wg�����6������qx	�.G��.}��=��`c�e�ZL�O��ܓR?�.w�@"��Qh����Q���Í��Yw���gKAt��6��
J�2W4ڤLIy�hÇ>v�N>�B>�7p�u�2p���&<���0N/sX�8�dl�!��A�-`��8%���x���/�!�h��ˌV�f�y5��c���``ǀ�C�c=��_^.~(���6�>	PB�"\�X�5�;������p�e��r9t�_^���t7n�e�B�#��Q��3 �q��$��t�����I�ʻ؁�.q��~��3rJkj���;����O
BkVA{ד?3�~T�m[�db�6��U�'�����a]-d8�Âkf�G�d+$V�Q�����Af@�D4��j�(cH��,�}e��?00y.�˳�'SÏdU�P�V	$����� Yx� /n���|[|�a��ɣ�h���%i1����#9�����ɇcwe���)��wݜ�)�{4�&�h�	�fd)m�K���7�p}���ۘE�5�Dk�ӝ{gF�6�{k�S$�����s��_��\�KI�D�R�<cW%��!"��ѷ����C�kM��׬aǐ�D���#�}5�<RG��_t8�������#�lqPN�|Fw-�Wz�t����8L��{�����i��w2����kTT�#�S;/�/`�J�؅?��W j�]:��LZ}[����X���f(l�,y&JK��N%ߺD�V^O�5��^o�6o�+�<y
�0��ַ�ɫ�J��:�x�*+҅�7י�]�~۽��{��ʎ���M��sZNWt��u_�oc¼�R��;���M��e����51]/���B���xX>�oЌ��]\�����I�.��Z��p���Ɍ+~sB���[�ZS�`��g��'�23�.�W�	�L�:��8���x�UA�-���
��
�V�����T��\��O�g���^��U��.�e���xT3{Ԑ��c�M֜�}�ip�W1Z{4�G{���2�����-���,u��A#�2�3}f�ۇ�n=���q�i���b#��B*��Oݱ�4)��vKjY���j��qħl��`*'�W�)>��w��=H��VO���}&d���v,�Y�j��+g�T�/��=!`���m"�g^%���j*g�Gw�1�o(]����R�<)|��J�Ξ�涣k7�����(mrK~�Uq�Q?uМ����
��*��E��9E��!���'���gv�1cP���6����g��v�u���~�l��DH���e�[� ��pٟ�'&&\A���	��7��}yyU�!Ls�&?�0#=$$wh��S_����p� q�� ���oU�OG��}�eh|^ac���%h������]�Ǧg��w�B.��yА�3���,����C���26@1i X���]�:�����s«� L��!	i�W@+��l����aj�q��\OX����mr�q5F��@�ە� #u�$&�/q�Є3:�A���a�I��`%��"�����uLk*�qSSJL/��x�xͧ�F�i_2@�]9��^h����p����#��E��F��&��Mw�!�X�;(�֨&�x�Vq�+R(�U������Kd@d�=�ŉ�����MC���q�e�n��z��� C�x��ލU�2QCfx�e�Ɨ׵9��,֌u�9-�:k,�i�rps}\n1$R�S̈}D7D��@����kq%�y�㬞��Ծm�X�pH�;O��L���p�T L/hcV#	�ߧ�*m�̾H|��@�N�ʧ�����hp�9$�KL��%���F�*��L0X`� |o+_��16GMOxV<"%� �t [2�x���_��!:'''��Y�
P�mg]aT�qX(H)�����^������{Q�o��2)x's��u/:<0J�IK%>Bs�L�%2��7�!��6	~���?��r�,+!�x��ZN�W1���L�B�kx����nX�U|
~�]�P�Љ��F(O�k�)�`�؛��j�l�K~����D��A�x3f�]���R6v�r�VC��vm1�u��-��^ �;���,���\l``��`�iwq[Z���R�$	I(�@˃CCC? $�9����+ݠ;�Kh�I�V��!1I�e��x,�}y�Z]��Ɛږ;駆�p��w� 	Mq���aE����w��ҨG�Xb̤djp>
�~ʨ�N���~Z1�6e��f�ޱ4�y����{���*�LC7Yb,�5�#Xo&H���븰D���h'`q�%8����2��l+9##�Y�]�6���u�@��/�En�A:T��Ʒ�p!Ȣ��ܢl�j!���ե\���8b��ea���E�m��R��$\o����_���� ��7�YI�J�N��$�W��M4-�iSp=�˅��n
�	rKQ��y�z��j�����f�/��r@�f��.�'HrF\){2��uŢd؁��sؽĒ��NFwf�|e���z�xЌ'�K$��B�����>����WJ�~h��i�c-
���I�5gެU(N��������
W����g�K��B_U�]���F��ש>��4�g��b���]¬�Ĭ��h���~�DI �� ��p�S�Hh�;|y���禯�JR�9$4i�\�!�\�x?>�hnNa�{|�Xo������r���O��B(>UK�qH�&���a���52>z�gr�I2H����k	�ח��+x d:����	������
�,K:_�r��L�-x2�Zz��O)�r�AX�&�;���X/�]@��!���Ր�*
4�X��������L�P:�pr ��䰦|qf���ъ�\.���gC�i`\ L>���K��p��:�/�D	�Ĝj�)���ˑ����������ɧT�׫����f6&c��+W�nC�@F�<ÏE@�-�vV�wNӑ.���_�Vg��l���X�KĊ�"��@�g��'���x���^�&	k�c�U�Zcϐ1��N8�׃���	�Y5/&s܉���Gm�/�ˁO`,"���w7��Trm�7�1��m^%FO8��7�1+U}i���Py���T��ɜ&C'K����>)�3��毟�P�a�}�U��R��H��;�?��C�0��x0�hO>&AY�q[�--E������ޥSm����f}���?~� �dn���K�9�������P��/Ep!��2�� ��PQc�Ayn�����L C�{�ӫ�n�:�O� )ܳ*l��p��R({7�	��Ҭ�������ȅ���?1t����8 [�5����w b���N���e����ٝU��
����~oeL�k 䌒h�i�]G';�����{��7l#�xJ�B�e��f-���kA���pN+�J'f��4���C�! #��"�D���ma�:Uy�Թ��zb����p�A0v�v�3ڂLVh�PWBx���MKq�\�[����=���s����^�皤e"�?��j��TꜪ�|��+��G������_CZ�Wgg�J����1 ]C&��O��G���bj��p� �9�/��OB��AHƽ���L;�=��z��˗/��ÕjZG�wɱ����h�qx;�K���A0�ղ8��L�[�fOO�Nfs_ܻ�D
���-���X�_=���@ZX�-�[�%��؜� Cc�Ȉ�l��t"���r�v�K��q���duN�Efյ�m����V��JjQ(J���H����!����O2���zUzD3��XQ&*�"�lR��UK_�/(���� ��X�aط�YG�K[ׅw��O�,�"� �E���䊧DI��bE�3�����7�7Y!� g�oS�z�"���#u�����J����f"����`3�zK[�&I�Lk�J2BQ�ۀ�Y�����,��s?��o;28������aH�4�}����Kh�jE�Jc+cZx=FH�����Bb/wat�zӏ����d��L���8Ѕ�z}�X���͇�.(�� W�y��q��`T�lY�����
�IԒo�3�a�0�����{��S��V�_Ǳ9�/��,B��v�6�2��x�MBy׷=�����	؄2�	!Sw͜1N����܄_,ÎU?>��4��`dsAE.�L�N���O�)��O�%=��=k�9%_r�哂�e��;��,x����,)sss�Uf�d����jU�UF��`@�����]�f����6���5�y#� �����+)�Rnܩ�����\���*�mS98���8�������dA��󤍡[��ҽ�
H�Lww�)�C@q8��(��d!�r�f��]{,�PN�M�q�_%���>}�̘�'M�>�!��D`c��q�i{��vG f~��
���	!|:ʄ�){�\ f��h&i��D�$"�N&�k(�*5�eI�A��m%�&Z�oƷ��/Q������3Y��kZ`��a�hY�����ǩ�%���m`�u��G�:;�x��hl]���f��ꂡ�����B�\v��|���9�m
 s���aLC�!l$n�Z�k ����j�2��b��3��	�ߕ{\��T�WA����Q�g>�.�=�Oa�\@;�j!�HS�h	V����'��%=�xn���4�,ib�@ �M^�[�}�˽�J��8�]��������	 ڀR����_��$+����U�ɤ^O��
O�Xx"=�ֈ�%r�[�M��j��ZB���r� R���61�:��a7:���D� oS"�˦G�}����%��'�؆�fUgF�m�y
��K~���X���+B�2�IW�f=�
���F<��H�6~��E[�|&���p�+�9��h�]p�?�C����[+.�	C�@�nA��Kr*VIǫ�$F���vK%>�ןΩ�1��?�kM������9I�t�������/� �i0�cF���[g��� �_�x����Hֳ7`Q]��YH?=�t�C՜��}UA��Ц�N�Hw������I��9��N.������X��u�Ƃ5n��`��&-��<����+��\�G��
E$�c.�e��㋚������w2���QQF�;_�:��b=ۉp$nB�n���bI�$�-޿K�����L|�N�'(֚���v�������V?�5��(Uժv���b�Ӯރ�ܡ'��B�{*i�jR4���+$r+�?@���N��������\���A�r�;=� ���hZ�-���&"Vz�����腓&���(�M�n`�\.@@d�2yYԣ��c�־��
e3���+R /~sl:��VȲ�}�{����rv�D�ba?��9����c�I���!�^�m������Y�}�~����	�4�Y�(�#�Q�1��!gvp���閌���'�m�RsMJ<I��}v�HJ4x�!�c�:.�?/��tLమ���?�_8��c�n��:�!����lNg��y�Q!Ό�#�����%��4�ϯ �V6-�~��g��FJī�j!bxօca���P�`���l��>{PNO�3��DBMc '_�d� ��8��?b҃������&���ύ뙋1���?����GD"��C�J�!jhy���b��{h�o�Yb2H�U%������Q�y�Q��p�+2�hl��Y�9������ݨV�0�pF�ǝ<� ��#�m)�0{䝔��v��4![A\���z�6���	��/��N5"�zt*\HM�p-o9-��\������ ΅	_=W�40���RɍB�7w�A`�t���JQZ��҇X؋S`��0��ӆE��/ɐ~���o� �eF�r�ɿ��k�ZhX[�l?N�b�	5Z��v��?@��*9�h���(�x��(81u_ !+º���J�h�����7Y� ���H�Q��J�$��^�=*�����\�W�  �몞�cy"� oP���W.�Pq��i���P09 ��v��$|�ގNJ��HҨ{T��~��"�f�I��Z��p��ć�M��x3s�H�����?5$�0ݟ�1�_�x�3���lh\��4�
었=j���0*'s��j��v���C���a_h�t1Tq�wzp/�t�U����X_6�2��r���o�C� ��>]���9�Ӓ��R"��Ȅ��E����HJ^��v=R��@��<�m�Қʻ��v!%��g�����%[/|��s���>��Jv�dh�ε���ĵ��&��'�?Qhz8*�|^�Gk �XHE0��E�BQ���?j��^%�D��|��}�_����Wټ'�W��5�y�䓫����o�-���p���_?�<� r�E���)�`q`u���1�8�PM�lG��H�C0��J��
@#�^v(P��"�����t��.C�b0\٥���{�^x�E樭�d~%$�*ʆ�1�o8�����	�待�FB������(��Lֳ���̅��eq���3��=*~
{��i��
 �I.74J¢�Ķ�}��*]�d�	9Iǂ1s"]�,��ג�Ǽ�J�2P�4�:h���o-4�־ѽ��i���1Z&d�7�;���.�=nZ�g7q��]U��F%!K��na
�ؖ���4p5Q��bΣ��e��χǱJZ"�s�.�"M�C����P%�k�xy������i�:򐢒�&�y�`��m,0��mM���o�-��b�5zZ�/H�ns��A�%������P�*c|?#N�3��G1=��Ȑpi{�l�c#���dRȝm���<���$��cmwUN{�CA{���U�X�wcB��|�A14�˭����Fp*$d�1�r3^��<�������gDu��WH,�}��]��}u>.�Y,��������s��fa�b������@�s\�>��ԩ�[�~_�A�q������4���jf�H3��[��"gY�K�ƟH�u��K��%�"�Kv@`���"뉜��R-2��yD&wSUd�Wd�,}���j�W�j6�N͎���G��8���5�x";�� }#<Z|8g6�L��{��ލId�^ͻO
hi8i߽���_�a�Ɯ�psf:�[�+2�4v�29�����m�։�V8a4�{&�W_k�7שN=]e0Z��Z�F���vR���O���y�����JB��$le�5��x%�P�����z�\��G���U"r��;�{@�����((�@\�Ap�v�&@
W�o������^�Z-����1i 5�����)CՅ�fm�|��%qr�c�]�Ľ����YtZ���<Т����� �@�:�T@����U�D��L�u��6ߞ&o�Љӏ��`>��HP�'�R�L�4����cp�tt���-��tP�1�8��ri�V�ҥt�'�q2�#�?0�
���B�I�= !='�]����{�r|<Y��_�蹦l�D~o+Aɖ�dZ�E\.X���'�U�o][`����w�*8/��>`�a�w��vj�ec:K;nO����O�^��%��	�g��΀���d��:�0����2��Pk�]��X/{4x�צ�]��й�\��W?�� �W�bvp�_zI�";kv��6�C� �B�������p(g�F��h���/��J�U1�����J��h�- ��[Λ�P(��Z����s�r���;r-2�-���	����t6ΞE�%Qyڻ�:**�G����	�����dm�e�ÿE�C���|>`��s�[��/3�輾PGEw���[��q�uutpO�N?H�]���E�S����ɖt��ыc�ٔm��)ؖUc3��OI������y<U��~��B�R�LE�S�DQ)���Ǎ�*$��
ɔ�c	J汤c<�y�=k�sNw������{�>����Y{���������{��诎,�jLU��	>O��͝D�B�}�}L�У��H�O��K�z�Xl�~���K�����؆O�M�R����.h"�~��+�t�H 
��#��?\1gH�B��
�v�	��8�V����T����.+D��W�v�H���]S������q�����A�e�4����؂�OH@�����ja��\Օ���>��D�f�s��e��9
��H�fS���x�I�(K�c��S)#��(c��3<�RP�t;d�ݦw�~Zm��p��P�L�V���c�!v�>������k2؅�y@!c�ߟ�ֻM*J�!���k>]?xG�$K����A�cZ+�A7��`��@bO4U ��|�^\�h�ƕ�I���un���q>G��##죜e.��~���q�uGvb�_�J����������X�腤#q�R�<==��� �	|��\8?�(Sr�Uׅ���C�g��{Ze���&�Un��>��eР#p݇1F��Z1�"i��)�p+ܚ�6�vni�kE}#P�X�BS'\ʶ
<��gP���Y�m���P�\�l-)7��{nB��j0	�����W7�d��\P�.""R�� C��{|��nT�M���l�ٽڢ���I'�Y	
���i�h^�ؑ酥Jߋ
y5FZ��Np_���8u���t�5�&"��*#�\jv0l�ĮU�kw[3�H���s=��Tm<a=�QQAS���ǋ��Qh��|X�߬���������U�ݕy��f�xC	>��؇hL��j9֐�n>� V&��!9����5׿�){g�&�dV29���X�^�����V[,�{��n)����X�)�U�5��t�ITo����m�[���s`J�&��F�z$�s��mj��::�v���Ô��nh{�f���[3�J�\�в�Ǐw�r������j�`�)�䉈��Hu�oE��Y&`�V��e+'Q�� ��a��xܟ�g]ݶ�\D=��y,/�-h������|���h��r��e?� YC�[�\�C�vb%���b�ׁR��N�w�$Wk��
�t��_�P:�u��� Uc�0�ᶰ�l�O��v�沾�5�P8�\{h@�Vq�F-�cbb"�, �k��
�ek�/��/Wc�tU����������kzǾK�LSZS���J�%�Ã�b��F��;���x�F�����Q����Bh���zbh�!�]������t�EH��E+	�[+����	�`C�t��D.g��Z.F�Q�8Z[��o�n�2�.�{/�A|��^�#ga�I��

�(�9���%�0V|{��T��z�D��_O�F�pd�ۑ$�ؠc�K��}�����@bJ�����\|e��]�����A�^�뼗"��1��������u�7�˿)�3�S��*�6jD��r�W�<�
���;c���=%Z�<���"qX_P$Ol(�M�>k�-�#ia�0��l���0F҄��%Rm�B��*Bw�f4�J&�i^�;�R��i�7+IU�a3<ʝ��"d�D�3h��&��±����M��s���ۀ)ڤ�9^��'�������e�=��76|b���*Ci����W�AO��=�߳��e�3,�vx;>�3���鼑g��G�?�}>|6@�1Ä0, ��J	n�M<���h��gAm��ryA�B\�0,!^�+��l��/!Hێ��<Ӭt�Xs�#�U�]�ᙅ
@u�T*z�a��8ĺ���Jx������f_����%Q�l_��M�,,u��f�bg�3���Sw,Pu��J2���Ų��?�b����M�a����d�\R6�+Gy��J��ZAsY`I�H�q�cn:�I<��|��w+�E]���<�~�8{?f�؇|^(��o�i�Q�����־[\��h���wg�ʥHi����7���9ԁ�[� ��Mc!1�{j9��!_��9;���,ļ�A�����(
�t/մ���ev!��b����ٝ�(:�iJ��o2��e ��c!z�l�]���V����R�æfH���IG��Dm[wY�	�H����EO놓�f(���l�-��v��,Um������C�4$}ꤌ�b�>���Ƃ��XO9��%���@�W!V���eQ��u^�4@g��1�@�a=C��``g¥l�MX�U�E��+k��:B>=
�����g�q�I�w���&$���X0�G$?�q�b�ޅ��i�-��28j�� ���$����| �́��5�Eb�(�:�}ؾ%����
Q65� �chF.�ŋ�oC���	r(��\��<ע��C���v<mE �j)�?�&��8H���	J�[�X��=i���P�]��w�0d�:��Lĕ�=������7�I?����
�Ny�s5ٮ*��AW���hP���2Ԓ�M#��T]�5WW
�^U���e
cn��F(�C��)�s�	h\ߧ�;�<�$;C�P�I�oͦ; �I�^>�|�᱇c���̡O;�
��Z/�h�����d]0q���G�G��L�)u�=YP ������[��{�g���z��X�]��$y�m��P�߭h���Y�U�t#z���f���e��;��\7�j��5�*�_M�(��[�$�T)g8k���*.��b6�"��^��:,�ZN���F�� $>���@q��5RK��gKw�@RC�/^����o2�������G��}M �J�� )��a�)��M�����ITfmD��I=������2����J���˳��}�ɶ��|�A]�t"U1��z���0��@���T�S����z=_{R�鱚�4�����;#�
�9A>�ѣ $���c��l!�O{����%0���-r�Pi��I���b� }���3q��!`��h��ᑑ�i��^�:�0�Զa��L��|��܄a�o��+�{0�;�E��b��$g<�w�S��e��L�L���:hՄ����M�ô)7vz��c��$LmZ)�2�F��|��,��SFn{9���(�A�{A�S<�.M;	�G0Y?;!�A�F��RKɁ}�ss92G	D3GVEA6�^���XIr��S,ĎH�����_�J�Q��ps`��u7��V
��u?�A��<�$���>���:�6�r��|II���b'g~'�0P�J�����p�����A�ډ	
��5U�E��gwm����Hܲ���mj�b�QzpF))�X��D��,$�xQ�>�/%u8O,�M��	}X"�}�����!]IHTE��I;��u_C�ڈ�{T �Vo�lC�X"[��Hq�K�jp����I�&d3C��I����z����1�޴�/5u�.�V�篠d5���4����{*��f`\-��̩}e��P,�Ӭ��jT99B�J���HC_sqNO�P�Px�=\T�����#�s�Ά	Yp+��S�L��J0V��H���q�,�����:@rn߼����+�[M}5Y�f�5�D3,���2��f/��Ր �>r�t ������BII��wP�� �Ky��E!�gx9(/�2�|�� �ěE�x�(�PN%�QN�:Μ�W!�,9�62C��,V�Qd
,�����_p�r�Iʯ�Z��#���|Oa��Ơcz��Ux[q�~9D�E�����*nSmc�c�ވbe�M�RJ�c`� ܨ@-�6��!a��M4�܄"�pC)`�� +\�#�{"��J��`��C1줪� %Y�w5>�"�s`��|F�Y=�`U�J�v��s��D�^�x�{�/��IQQ���s�9�"ŭ̥hBkV	�@�fv�w ���-b���WQo����:8Iυ^C�9i.��?!X������ÕJ�V>��HsqW9T(��:����.��%�0\��>�Ts>���6T3�hZEp�Wx:�x���cG$}��b<>:��GK��.񣾞�O�8��V�N��HJ�_�^����<)buސ�!p��Iw�3(����Y�B� JI�C�9M@Up鉭%[���e����Ao!I%��ډ7բ,"�>R;�I(�r��W�������s��)hIBVb�ɢl��#74����}�Y���D��jj���5��WcU�U��TT��9�p�MX����.Fj�P�}��l�����e����'PAck�H5F���8���舢U��O��Z���Pt7FM����q�M�R��}t/��6ˢ��M�b3���p)�xs�����t'Z�g��@l�(�hM߶���znL�b�麅�S��������#�2e�0i�L�&<*RW�����NM�UXq]��R<��ϔ���&�;>M�)h�K��c���Y+�8��Cl���.Q�`�xG��\F
f�4�]%7����L����˛��چ��N���UG kB�*������2���Xj�v|-���ީ�w>K�@��H|�2��1́o��Q����m?�s��nBxz�|��|��b理5k�a��[pSs�����#8�A�'7�t6�=Z/(����M`T����z�ގ$9B2$�Am����)o�ȱ%�a�ނ���M�%���1jU�.s�@��F�&�� ����1��|Jb=�0����A)Z8�
�k֨
�P�ƶ�"9Z�f��T��\�T ��0�M�be.V�R�.
��rz�%8A���C�WX�Z�WJ�P$Bqkv�	��5d��|BoB(�2��N!�HL̡*�����!{��H~�G�C?��pގ�,9��	_��V^M���n�8!���@��3��j N�t�`�'P>�TY�Pi�޲>�̈́�m�0�d��"yxA�44�YF�}7��wʺ��. ���~C6`��<
@b�.Y�W\�̡NFD��j��x��g+�zPF���	Q��ԙ�0�f�HS{%�\�E(VE(c�R�s�~(�\r�����+��O���9���T����Ji0X3����$i���@�"����GsHWX[�B5Zoۆ]7�\�$�Yyz�{to�������*	��x����"u�����C���aX�V���PMa��Bf�cᕷۉb(&|"��|� ;�cMD�ɵ��7���#5:ٚK!��1֨m�1�y�C�Л@E�/ �;���#M4��3�S�&dG�HM����qZ��{4��܃z||�w��Թ��z�I�Gb���o8�(��2q<L�s��c�����̫ E���"՘��^
�P	��赇ˇ������/��G��#v��ǃ/�o������xmZL�P�#��ky���3�j* ����ԃ��Tc���E��k�W|e}]k�E�e�4#�M�B*��H��O�Me E!��ԸXsg_l_� 2F�n"	��Jȫ�65>�ʀ�h����o�%��4�N~��ޢ:�n�h�P�����s���w ��WJQ�Ձ$��JGٌ���<��� �7�a͜������A��X=S�n� ��x��s��c��[�sC�ч���>����V%Si>(xΎ'^��*��(�ؾ�qtޤ���:���y��7A6�Gq�N�"�ɯYnή_�)�FC�6>k��U��+
��Zl|����U����ʐ#6��L ��Ύ��cZ�K���"i��ƍ���!��gkW�����M 1�^��n��m��z��V��56�mH��l�Y�w��6=�����Xߛ������-��y N�q�w:������X�P �v��#4Ҿϻ�k|^��S$��2��7(s�F�8?��d����A7P]T\E�-���g����2Hӆ:��5-��CS�B��W챬����צI=�u�s5!�����{�2�`��̲l��+�A4}�?+A�k��)d~�����v@��c�S�G����MWs���d���~_��eÁ����F0��kf�vr[�Ү'_��}u��������{ʴӐ����Ⱦ��k��?�X���
Y�KF�<2�Z#��u+����ւ;�m�����u����@��HSEČ@�.�و�\�?�3��h����н��U�?*e*�"�:/��,O�^M ��r�&�Q_�'n\{�O_b���bv7���#J5FHa����Ѱ�����Ԁ�&o�|�*���n=�܎�3�D	�G�������~�ߏ��~$�Tu(���8D�-�OmZ}ZcO��⺇t��8��"�OQM󋟌MU����h���X����]=zϘ���4~�?�u��ٛ{�����M<��hQ��%�U�Q��pt�ӾضsDj�#Ƶ�_�!��gb���+�*��wq�l�����]7���^���������]��K�?si�i��˧�������ePr�ˎ�X�KHNNVB�Y��W��P�h�0k����Ǩ�*�&JYu�F:�OՏN^W�T�bR���i�_F���C����U"�Ý.��o�R��o��,F��<59�>88�pN(��1���(��7�y�{ү����b/����ܻwϽ��C�;C<뺁��M9αƞ<y����´L����j�&����&���G]\\�ǀF[h�������0p�jp�t���je�Y���9���%E!jq����h?�H�Ύv�V�_<������纵k׺gx�,{��Nu�J�;R&����>n%-/�E��¯���P��w��o˼]u{������Jzzz7��f�n߾=�ۗ���o�98$M��uݾyS�z�ȯ�+�ʦ�~Qu�P��PTM�ի��z۬���c����n�9M�V~aȻ�[qʯ!����r�)����J��1�@�^��]����7�Z.�u������v����٠
���և�e�D���	=�{��y(+j&���ye�|���c�jWW��ٲ�h��jv�o�d�R�D�Z��!w,X`n3=I��膍����e^)���K����hR>���͝�����[�edh�)�`^�;�{���ܖei(c?�5�P�A���i����j9�p��h��4�7��$��������]>h��)��7���r��`����L*Ev���7b��e �ˮ??�u���c��0=��<J��kK�y���;Ff'��8���;��J>���/�n��u�K:�\%�T���V~�E��Ƥغ��n���aq�Q�量+1�"#���f�>�����
��m���s��Ϛ2�p���b��c��)������C���
��s�g���Mz�f�����v��H��)��8+�����#��Z����22.5���z"!�eee��UW��kփK3]�t_�"##=$�gc븽G�߇zzz�<S����S �'Qko�i�� ��o>+&	Z��v,{α��SVV��E7�<;;��B`��Q]f��t�;��������xw����2ه4�!�+�
�(���T�hh�<������	---3#]
[s�k����k��������Mj��#�@��`��촴���X1hD`�!�[�ܗ�Ә�EˆGM�K��ι��IۡX�*ܫ��iCGG��f�&�fv����˗/7�/��Ɏ�����>�k��]=Š`��p�ެ�'���'��+o2�[G�}�����L����{{�<��^���Xl�e��2ao��������G��E��JQHH���������p�J��ğ��K���t� P���'jZ�M<��|��m�7���&�QU��: ���Xؘni�u�Б#S�?~�������ӨE����8T4k�u�֒X��Pd�V@�d�-��hg]��Rs�Qy����G^���`����@���הEB\���e����=O8th"�"P�<�͡U��\�����S~���ﲲ,�Y�,uy�**ZQbbƈi��ĎvHF�����69�s��8�U�h�Y<".&6� � ӋLP��k���k7y����RXX(��³h�Ql4�mB��]�����d��ڙ�[2�۫��D;�<V�������9W�v�����.8:� �t%��WɹL�r`u �.!�p4x�l.��Fw�������J�9���W=:���/5�Bwz����`:ˑ�<G1;&?#��8 ��mxg8�~t+����L����Ǟ/����mg>s�l��x�<�Uo�os�C����C�l���)0��Ç�W���gQB�JQ=�G �M+,��6ض޻#F/����e��\歙 �u�� dT�#��7lX���#���oL�S=v��!�0��K�Di������|���煃U\�xLO6�ʰ�v�*��T,0J�n���=�W���i�egg'g�1S�<��K<\\���AXZU|��GEna6_�}ripp�iuu��>����ѡIo�=��������障�Q��#�%iu%7%ed�t\�5�SB��ϫ��.���c��Q�c���'�w���FejldddГ�\��B�YqF��c�������]_�%�<�O��HH�m���|���I�\���KGr��]`�j����7o�p1y�D�MG�e`�"GKmdf^���s������Xڱ�no�!V���GTw�h���r!�e=q.(��s�(���E�'&�w~����xl�8j��ó�WSSӆ!|�M�wt�~�����LLL(�����~Ѣ��N-HU3h���pp?�/"��T�;#J����@.�<ݯ�Fq	4�RRo��y+]u�c��|=�Eb���,���ڦ/-/-X�(<���T���c^����vL�9����� .�@�1arp� �1vƼn�e|�귺O��x�j�d頗ͽ��k��8�z��)�oV���ǼsNZZ�ѷ��~�ɣae��+�?�o���o`�����M �	d�U���3[[�Z����3���(e��ny{�ܞc;B$�XV1?0MN���PoJ���=:�Ou��)jX�x���xRr���S��mFV�6Rnab�7F�{�d$J�i���T�xo�zmr�B��Hs����1.�rVg���1H�ēv����,��C��=z��FGG�@x����\U!�y�0��q��Mr��	8��Z����^�EǼs��Pe�)��O(XH0�����#e�k"dt���_"�y��x `	/v�b��))�SM�tMm-���ٱh����u@� �C�Qy�� �ۏ�3�����8���71,y�����yh�ܗ��׆��xO???s�^��Ml}��h�d�]�H����l{2���^d�R�:�3��Hn驩V��Ư�4����"����-� �ج�kןx����Ex���o%>#��=�3\fȱ k��1�R{<��`��<�WYY�\���>�ݻI�V�.�-VKRT=�P+wssS�����x����Gx����X"�|����b�$��$���v}�������	Z����{0V�s��e��U	d��|�1��/J�a:&{o,��@�E$d��4!g��y��V ���y����۱�222�A�T���Ŭ8@A q���@�34��w=�I.�W��n9��q�<t=Tm�"�Κ"!z��S�����':�tXǭ!�޽���#+�KeJ��'�G�<G�XqA0/�́�Y�<G��H2����r갧�'��Ĥ����z��#����@<���� ����N�/C)f���" ��Jq�g��メ(�d������Vb�' �(��Ub���2�J���ۻwo!T��<��
��[���y1Ӳ�}xB�L�&�xoN	�|'P�+G�Ubq��C[����Qtӽ|�;*/^�ݩ� ����qȎ���}}E�b4&H!R�u
�=�s�'bLٝ��zm�!�� �O���qZj'j��䏲��O�I�T�{��3Ӽe��S衮���]:Ve��[j�
Y����@SR���	�"Y@ˮ�][�Ӿm�� �.�y�իWk%@z�&x�2)i�T�ә�۠�f���g$�tKU`�Ť���ֈjcЪ:}lх�#~J1u�����mPw-� �0�}�Mu
kT�R�Y�\h��E�u�@#V]<:�Yut;x�)��ι����X3��YOp#)����ў�/_&_HlC�V���[��Y��!�r�ܺz�ƍr^�Q�`��.��3����Ʀ���-CiJ1�2vLu�?I$Y�TQ�-?&�� !��@%y�(ݲ�p9�����}���PpΚ	����Z���\&{��kAJ��}ll,뻤�+D-N�<�w�ӓ���1��o�~v�ٓ	Z�[�x���	_�����`6`�4�r�a�<@𛾀�]x�]�.1����յ�T���Qǧ����ʹ�ndԣ�K#|ie���ӧӐ�<��nC�����Y����u
�لKI�@'?�����pI�"Us,��IU�/��0��o��4X��
��n1�D
�#V����0���|g�Ԙgn��Qf^�řr��>��Ǔ�L��ױZ	�f;� G�%D�p�q:�,Hluᐆ��333�����A�VY
�t����h��x^�L4���3����P�Ǩ�K��Zv�_*��NNq���x7s�!@��Y��%��:Յ���"��}��)\�	�h���a�uh�5���i��f��5;a�`ٵ�9�1�N��״��H$?���9矟B����^x@U݂���wɚ+������ӧI���:9�J(���
'W�Å�:����Әx�A�h��}��i�1�������~�����_�Y�.!v�Uf�}�V������d���� dO7��:͎~C4��h(_A�ӧl�;>|���j��!Ë�*���Y��7o��p6C��{&%@h��@��z]�K`CI��?��$%%m���6?5�lٙ?g��E��p�a��I�G����)ÞK�}���[./''GƎaSH,�p�O���8��Y��!��s�,J�{%�PQ�Wh2B��@��l �IOCB���c���dd��jBO��w�t��3�q�^�ڕ�Pub!��d]��А�(��������4�S�>�t,O�{.���̔�u��̂4�fU��Ie啃^L�}�T��8�F�T�� �n]up�.��Q�'X�����Ւa�d�r��|�BO�²1�">���`��Ƣ��q���O�*�^{��`Z@]����?��sƕ���"�����`B�}0KB8��2\S|��Ĕ��m��K �Q�E���J�}���*q�F��nEPT����Cpzh����;�R,ѽt�5��w-�,��i�#o�t��Z#Tn��� Y{k�â�L�|(�)j�xTΝ;���S��ꬥ�X��������&
�<+K�Ss!Ե�������a��pLB}�^Ksډ�Aĸs��*��U�4�?���5��m�ʴ;]���󈄄�^�����b�XO��7�=���>x{�	�F���[z'�jA�������9�>b�o�=��n�b�U
©�Gr�C�t3��pJ��p�( ������J
qm�/��Tz�Pqkkk$���&)�;�~��Fvd�����A-h��\^*�>�7�yeif��ƍ^'|��˘_�����H\\\ d��1.%$5�ne�n����3Š`@�?����c Z��.���2R �������0__�q�K{{{��O��EF"�=����{&��3�$-!T�;I���&�?|�(X������^��t|yߠx�e�Ͱ礝�� #a��djj*if��C�����S�ez�E�ҥ� �c9�d?���b<�:xZ�;?>��M�A{ɪE&��jj;:���/�̸4���ÞIzYjQ2�d����;��hW��L eY� �;_�����]K��!�wbN��ؘʈٳ`Y� �P�����*���;??��2��������}��˘�z@��V���/�t*.5����aO9 i.���5�رc����ې k/p�r�uk�����v�*#�k��W)�����k i�			=`}��Λ�w�a�߱�A}����*�"��i�u�3,*ߗZ����J��y��`���^# ��)�9hpS�J��pZ��|sf��\\�ӝ.�H)}�������EX}��t�UUUh��69�F����}��90n?s���da����#h�Q܎髒|���lO@���1�wGa���˗/� ��%pR2]}��!C��[��8Հ�l��"U����ðv�{]}��(t�h�	���]�^�����Ӄ
��4��R��r��nk�,�9@Ƞu�!��N|~Z�]�u����R<���ۄ�'���1V>!���}�L���w�����K�7�-�ɍ*��P��T�v�^���R���r҈����{�%4��E3̞���(��MɗexO���qr�oh\�ʓe�������`���i������u�[�QSu��>r�Mo��*�>bڒ�8pl(�v������C&P�"�٣$H��c���L Ä�{&A�����	��*�����R
��&���B@�h���]���Py�;��Q��Xc���%>,�]>|�U�x���_��"������
�� �B��~���&U{m����s���}||VD'C�^ e�G~~��&�u�%e[�Q����J�����Zu7���~������m!��z��#E+��B�6(���C�IR��V��[WAȡ�� k� H��22n�e�5��/_4��V�_bEkjj"��$Yi#$�n]��&)A4j�Zʲ�ZV����y�@ᮡ��/8A}����I�1�}� ���Zl%�X����FX�@�Nk�x����B�^�vP�8���M��F���e�.��)?�=gBK!y�K�W�ሶة#;s�l�>6��OȨol̔�z3	���4p�4�V�"&]$�}0{�~B�ID�'<2R�R�V�����FzK���f�C����p0��|E W'�U�C��#G�H�&�P�Y�_�����O������)��>F���?�#0�[� K�ד{�>ntt���Z]��]�F<8]��(z[ \$jaa1��"�% TP3���kkGB�ސN���/��)�]�
ɦ������@��*�:��6Te=�%�(��a�%�=V԰�U�n�F�.)���7lX����׾���GKX�.&hIS���k�*�������	��a��ӷ2?Nz�)�vC322D���1�����n��ǃ(ϣ}�������".����� ����H?��,����*g��G6�����/���p�����-3jt�h�c�1h���X���K���I?N���a/�*�ہ��3��sn���[ɾ"s?�G�鑳mvyc��`ڞ��Q�=�Wֽ���g�Pr�|:���kF�Ɋ�*�n��*���Bz����{�y�`�.--E�����K�H;�(~��K�+I�j�1�疙v i��*�>��e �c?~��[ �^�푔:t(���f���Y0Hc#/�7�>�+nz���QϞ͞p��VR����V�Q�7���x����q3����q��g���"!����
��JrpK]�XM�%PtK7Q�yí�L+���󰰔i0�;�S�IY���@�qǰ/ә�`����0��6��GY�LȦ�c9��
�a���~ժ�����;P�)�z�
+�)��P�~04�SmmV7�Y�]`��`bb2��[��U�r��iZB���k�����ڳ�@��=v�d��ͭK5V�q�|��Ғ!�V��
\]�2$���..�N է���a�&w�ܩ��@*�1�S�"�gH�� q?�k�`�m�N~C�͵Cy��3��Y�_A6��Oqh�<ZKHۛL�3<�x�����$����\&�9ϟ?�+((����I��T�cǎ��������<R��>QѦ���, -�U������\�3>�9�;�i�eC�v�8=��tD���@���NW�!T�ǕC�	��~P(�(�����������N�: '��6q��y��e ;!C���Ψkh��IK��c�� j����ɩ=Op��c�r%���ƾ��G�W�)�
�A��o߾ՂM?쀄��Uei�Kp������#G���H5�������Beb�!�Z^Z�C��}),,��GS���xlI5q`���.�N��N��?�8� ��`��H!;L�*Ctw�I5�%�(���k�	sgA��V)���6ʳldm��`.1 u��x����Ւ�{�2^M���^��3���LM�nD	 ���+�:5vw/��l�*���s��M�k`�<)�M)Q�6.0�}�6?�b�t�9����82�un|�Z�.'&�)�/�������p�y�LzL��ń��,h\��l�'�ړ�ݷ������ݻ��J��QQ㧰b����Y���4T��kiӭfQ���A_K7�-�vY�
o 0�b(oo�yOOO�sہ<��/�>��"#%u���^;BX9H�y��������Gt�N!�F�M��B��&G�,��`/\�_q�v���/\�p���< ||E~��1::�~L�`f�抃�ە|9o�����n�&P�� �B�WU��%�7"(�����O��6�?}�����v��H���J��Rrr�""##y}�D���~>,�d���}ڔ���q
R=]�O�`\˾��50ۍm��}P�D�W\]�Q��K/5X���V\_���
v��ʒ����j �j��
�x�!,�j Ԥa�Ȁ��uu��h�蕦ࠃx���-�S��5���L����[�#G���!=���+¯��� �
�bS%�i�;	Tj�ּQ���J#�0�q��pGggghB%
��ADMS��N��@�#��(ds��4���C�8����j|�����t�������MT^B3�q�f���+�p���orjۊ������)�v�q��C#��|��h�7o���1�E����2F����q�~zf�/Z��03E�;��&?�����o�7b�w�V�CM"�o�^�v[uR
���_�"�3�z��kkVF�R_]̱ofO�g��w�+��S ���ˮS�y���\��)O�p=3���r������R���		.�Cs3���n@��dKNɢ��\9�i�i�Q&��{�Ϧ�U_D'��AiB�2V��RٓgϞ=���A:�>���Xȃr8�W��:�'|&''��~���R{�y�@9Yx��y1�j����[,>%����~"+A�5+�n' �03;�� �����y���II��s��z{�x\m�rjQ|M���G�._�C�^�}���@P�*H:T�GO8=~��ϑ�LUrs[��,�+��}A�s�m�im7?7���e�^uu�-��-��ݓF��@g	�O���T�����젆� L^�~�G�Z�/�jԅ��GP����_��v�b��!Dۨ[fff�o�^-t����0�\я�C��5�N���n�����B�6�1���;�������Z7� -$�K�L+V��߾�$�8�ف�x9�okF3�A������g{�T^����n�́qJ1��ոl�b���D%�41II'�_�=B�"�;��*D���]Eq�ۖ�D�?�Q�T�_MS��;::V�w�R�0NOa]���h�ny�!a��K}��>6���J�t����%�ʩP�����p��*?�7p��˗/����!;�k�9�#G�a)q��J�}���1h����q��iG�-���E�Ղ6hμ��~��cqqq��]��S�琉
;�����eC������ ��>s�-q�v�=@�O$HF�����B�N'Y��䤝%޴�����d�psZ�KԴ)����s�|$�R�}����:�nq���@��W::�V]���PFVV��i< \e�T���� >���ۨ����S����꾀�----���Ǡ��v G��xRN�,/�,��?gΜ���q�7
�BM8i����-�;���XF���Cg0m ����_��qs���J�!w�\z���s�U$ �e����c��O���]3������I"Eq �f�����Eź�M??�� �}�*1����Pz��9!ʋ:\��,8�r����U�ג����Ԉo~200P���R��6��QI��W��MN��_>�<v��B��ɒ�/��hB�=>f�>�;��QB���ԏOL�K�
�T@�L�`}��H��vmmm&H] eu7�l=��TT��q�v*T���z�_�����$���zB5G��	at��m��1�I��ހW�^�+�M�Ӛ^:�/�ͤ6�a����ܶ�[+�D�+�|����g��ݻw�^�»|����ԓ������m:���C�Ӵ�F�:�R�TfFVʍ��/C}|@\|���!��YXx/������B:�weW���BeaYf=�5mp��f ������o B/�T2�wH:*���q�����}	2��+�䮢��/��$P׃x֖�ar=UFΜc-E�abb�yOb���o����4�X���W���Z*3��V@��[�Z���>F����J��|T�q�h�M�S�k>*E�^mhl�&��rs��K���
�]"���K����Q!|r�[Qz�D���|/�LW���<8�b��Eo�!�SM[��KK������>#E��8���Ń�Ν�iCx`�`v�!��!>�Бwi;�Whc�|�ܷ���޽;���]��(5uuG��'AW����T\O+(X�nll4�{Mރ���}�`����w0�`����zĨ���v��Չұ��]_����������w=ހ����&g�2��*CtF��r�]ži<�G��T��tR�z�t0�[y��Pa��7:TؼQ�t�%:�������uuuU���ZS���Bt��GoUH-;U�#��T12ꩆ����� ���lڈ��43R��+�?yrrr�6 � Ȫ_Y6l�ϥ	��4����ӓi �w�I� �\�{�k��,>=�=�1��m��K	G��
��
p���3�	%E�~;����A���)U��Ă����F��,�1!��
���軪�\�v���)j�oe���q��JG;;�f(�� ��z�>ԋ!P�S|�:`Y�s����IU�*-�3}�E�ݍ���S��i-by����ec�UrЮ�":
�s��Z��3G�� [W(>p8"v>|��ԑ#S�8lü9)�p���>��#��$iǨ�aj�I���5ƴ�5�z^}id�%���1��3P�	�?��W��Cuƻw�C�����T�ct���&.�������ԑ�4������"����:+u;���l^$ltuE�U(��z�����a���P ��;��H�ٯ�OTD�g�<����r�Ǘ�r~�������6%9����h����drS}�h� �;wޛS��ß?�"L�T�׾�O���4��G�؁C�CV����-��x4v���Pg�Ry��A����#�psS�A#SKhj�=ǖ���d�_�-�2u�t���Pe=1wȤ&=0 ix��&6vv�{�X�Ԧ��T�������˗� ̎ ����6���� }%�s:lP�|��O!�`moJ�{����@���J�'=�"^��ᬕ䎼�n"dJKP&7���H�J$y��P|�H�\-aQ��6��<���A��z�O����q�6��Bm��D:j�e�!}X�A�?�άm��ha���q-lhn�m��0���9T�����r�z�gX@���
�}���_`L��[L{گxD��pe��X|�&�q��v��b5��/�UPc�+!9��EJʈ�\ �#22?�,��
��pٝ���z�Z_tg�NH�ikk[p���RA�_\\܊����}��C��Ǡ�07���}"��Tg��Qd�Ӑ��LLHY@�l(P�Z�x�[������yiS^����h���:&!����Y�uӞ���Ԟ-�X�¥�2�ֺ�P��~�_y���kH�T��b�j9��F?	=��=����i;��]��x$+#����͉sA��wX�(�L���c�Ow������g!�(�|V���,��To���ӌʓ���:7n�*.�W���Ϲ̐����6�y�9�s$������H)B�J���-�[�ѮԀ�;ck;�W+7Ӯ�
'$h�ss/��*��� ����t��}~;���	��A�2Ys�̠C�{��(Zg���G'�@KH{=��Ϟ5K��.^�*�ƃ$��6�h*>!�A���<���/4��� �M�͝7�@lhhF �J��R1��6��J���n�,��(�2ɉ�	��̅���q�Sũ�*��!�\n*pE���>syyy���ʩ&�
��o뉘� �W͹���������[��m���~��� O"W�in�Uq�m3-Cð����)���Q8y���V�������������ZI�c�&iq�줤a^fn�I��M#�0����܉6�UIII+�Y�*TB�]�v���a_Z�lx��oL���UP�(F���`H#�� E*�8�k"dj#dfRPw�||jϞ9�x��5x����{�22\����qD+�X���)��/����[��f+�DBq7��+S+���#c��<s�r�(��3{1���ӓ$/�'�22��'��_�A	Jty	��&D�G�4���F
Y�!@̢�w��]{�Ķ6���Lqv��С����;�@��.Q�r3���� DB w���Yj!51��=�*7�ח���rPG�$�߿@^u�`����}^,����A�S��+3�(*���A�Nb�ܱ��f�����k{��(J�{*�*os޽��?�M�J�-y�\<�� v��v��m�\��
��g�����yPCT���-x�8W���J���Z�$�E������֗a��2��'ҟAm��ǩ��$���u=�G:ȸd5�G��"�*K6���-�z�W�NTK�B�i� ��>U����Dn<��J8(��RH�\�92<����(���&��Z����me�󅁔�$:J���{+� e��-"6��Ξ/))����2j�}[�ߒ����?E���J��1j�˞��.J�@�zfӧO�)�jFi-E�����o9�$�j��Q�]����i�/QR�?3�e\A�Vf��j�������`N[�0�z&}�m�����(�Wg|nџ�Z��:��H]�d�ޚ#��S����c�>j�3���/q{e����݈���MI�u�bbii�]��Bs;-z�;\Vz�&�g�L�����������[�Z����0������J���Nc�2�k��#T�ji ���$�]��	Ǒ��u�Th��|�Z@<v�X���磨�e��<������&%��$�M�+�T�8�x�а�Q3AK2��7��4qq��ׯ����n�U�AD���cJ\�5��(?�
���!_����z��U����eō7��]��������=1&�.����倔�8ˌ*P��kkkW��j�R]S#2�΃�k��m��i5*��%ǆ���]٢���M�'��2`�6�9��<��³����`ͯ��Qa*yձ*Yv�ӡ�� �Jm`E��Z�#����WI�����؟���t1q��$M�C�e||<�ҭ!5:��;A�!i��
�YT/��!��S���G&�?��1���l���~-�����<���n�fݨ w����Q����U�<����1�q�z{���}GN�
���U�u�P�0{P����B[=�6ll���(.��Aꈭh�[-�>5�WM&���� ��@=?E]��˲�����̋�_4B�^۔��&Q��TFG��	oI��5Xq��)_W0�	 S�@FB)�?[d��=������ъM��Ѱ�y���G�� e�WT���B9�ҥK�P��&&Q�P�ւyr�qk0S[W���)zzz
�FEy\��uM�5g�b��Ke��� S3�<n�Օ <��U^`}�+=�ߨԣw���q�Ň��Y����`3���j(C������������/�q��ߎs�A��R:�DR�䄢TG��$���ގ�hD�f��4��aG*%�������n��g������|���Ϻ׺ֵ�u?Se� z̲��}M
(^�'�|�
/�έO�����G�0:����Jv�m
���G� �8�C�ƈLU5��TyZ�9��oܿ:�I� ���[[[�n��?�/z��%���Q˂n+3=�����(VU�<,M:��������R����]��ON���%h�"$4]-9=}�/ee������B�F�9y�ض���Q�?���H�Y1�����5�+?��Ĥ��_��]�a��齷��}�(c�m�������ق;���(���T�BU$���� kgi�I*5L�{f��E��弄NA�WVΎ�ܖϨ�9��r��m�!U�T`Z����|�:g����T___���{��%j^5�*�E�f������?�뢱�_�����ϛ:��m��?<��O��o��y�m�c�D�_�w=rR,�HHi�����M���{��3��A-��%�c����G��0i
�u�ɽ�����}�|o;�F�s.�Q�|2T#Q�6"�.q��u/���hH�nlè�Ud	��N�	�s�.������K�-������l�k��~�A�m��[�Tv	�T����{�*��1/��������Cw���qɛ�A^si�D{�����ĺUw��(��'P_�zl�wvGX5 ��N�	�0욷�Ֆ��%��S��#�9�.���y�a��ԃ�r��u']���\��_��B.m���<P���i�xG�1%啂��T�Kn��=��n8�m/��Ү#o����%��ܮ��������F��,�s�o/+�>����/6�Nr�[�4�j��d��J��|"*s1[O!�	<�p��N|^c���|qJJ~3Pn�"���|{���W�>�	�� �IA���-��o�����7ӽ�dg�;��x�7ǳI6�ְ������G/t�ڬ���? ��ؠ��Mع��I�ؑ[[VS������5$�[��h��u%cn��=�+y���D�e��Ӆ�i�rB=a�8'�����DcC`g����?}n\�N�/�S���nw����S�����f
f�/d�]�Q���9a��8k~�5�����8�qiiY�����zztU�>���r2�x�T|cK�sA�܂Cu��Z��ʜ�.��:yeq1|��X�s�y�f�B,�*�/xTTTt݂4ؼqf�����aݖ�{C�T}� 1Ϫ�zt����2{ɠ�����>�e����Pp:u��0�1?;<l��!��6��L��.C]��'�7�k@�Z��z�M���vN»▄���ƃ'n�{c�K+���3��T^����Ymfk;l4���2IK:���Z�F���y���ύp�`�	�ps��ԥ%�]
s]��=��Y��Q�K�H���kii)�J����u��������e�e<�|cC҈����}d��ٳ�ڟ�N��7s�J*��J�JeZf����K������Ӧ�4�������KO�; Ȥ��8��+���[��OM����1d��[ތ�s�Z9zi��f��'N86H��av����{|�X>?'D�؇�g��z�P4��';�^�JL�w6d.?~K4@)a������/�`��,��	5��}�
�9�E�Y&���z"=DB�q�ev
���W�wŬ�y�Vf�M��o���;��4_��x��4#�6������j �3����7�p;�
�dM��V�=�����F���3;<��@���X�N��3����x�r.�	�"�j��WS7H������Z���>�[Z�L��=��~g���y�XDi:F��+U���l��纍��ɦRxT�M�#.c_��e:�S���AV]�P�V��]�r��~x�%EWD�qaa�e��>Q5�$�}�Z��<�?������8=$�����S�C��ts@+%�〖�&ݽ�"�KK��q�=�KA�����J�2�Z�ޑ�l��g^�n�mh���4�����q����Ǹn�&	C>��ի��Qi�k�IIIi�E3�*M����L+��5$���_�vU���k���zA���ck�|��h`U�0�m����fl�]�m߿;�C'˥����𷨩��b����#Lq5~�ܭ����2K!\�y͎1k�W_ÈY�~���V[KK���F�c�;cccG���_#V�Ha�n-	e��yכw�����zA,��b�:�V"ݖq�ۻDu����ļNK�Â��BJ�w�5�M���c��Y[sm5�ܾ����Y�[̯/�gX-*	=S��k5L�ŹС��5�ѩ�/����G:PU��eUB�f�^�5�R�M�"p�콋x"Č�s��f�8/XJ�[_��&Vc���	x�<bF��H��i\D��0�9p3���35�o\�κh�b	�h�>�x���Bh���b�22X|+�8��Bv�UO%�gM/��;|n�\��x�*1�[rFFK[[[�I)*I�y��*�����/0�M!=olq�|RaN��v(u02������ �N	z��>���엓�佦�������|��N�<�P������?}:�
�~nf2�����:��i�Hmt~��������k���o�ߠWh�qWO.}�hM��ː���h�p��ɞ�Q1㒢��ؚ',HҮSixZ��J 0Ay�`����W#�(ZM�t#Gj�4H�8Y�~�k�F����������F�'�8J�o%VJٴ5��#ص�X
��u�#6�ZJE��+>o|�}wu�hoM�p1����?�sƉ���W���7uu����3RR6�bb��|���F��H v>Gj�����
z6)m�~��ُ�	��Q�� ��I�f���y@�	?���0K�5X@�@aC�Axtc2N�y�{���Q����K ��B2��Nr�CCC�x�m�}z�;w���rw�P�(���#B�mm���W㫿@��~�Ğs�a?'7�vpp0����Q#<&���&b�i�S���_!�	���)o ����ߎ��G䈾c��,�I^5R�F����@�Z����)2K���՛�7��s���z�,� ���<��۪ �"7��W��0�Ar$��]��I^��{�C�s^�2ؚ�/���1��(��|�jg���}xn� B�Ϳ���]�B����Z|w|RxD�� ��Sa;z�^��8��E���|�Iȑ��/ �9��]��!� ��>�Yzy�z�\B�#��z�M�rvO��I]S��1+[�L���fϿđ-T$�����Y�� Ω���c#ȱ�c�{M����p
��:�����c�q�y��O�^�ih��MM w� F��E�&m"�n��o�MMM�ڶm[5�IMMM�W�\yB �����oNwJ�tP�rY%^��q�l�MN��^�b�;}��qr�]���y�8@�%�-�6�ܣG�1��h�c�4���ȳsTe=*y��� y/ Ȇ�S��NȒ�₧O�8�"��_�� 0��(�H�B����N#�וؤ�o���5��["�a�����zO�X�آx奄'�����uP��KֈO����N��{\��&���L4%p褰F\�r!We�ٗ-\\��&�@���V�?���?a���@�C�ù�7�%�)�
O����5׉���#O�43s��@���l<T�"�5������<Zz;26�]�0*�w�7��rԓ(�v�*+�탦	qY��.dGӱ��	uJ	'������� �!V����Ɣ����)6���c�(��m輰�)����zAWCpds����;�1ʤ��4�䎂�\�������p6��r|8�����oB�u�4�c��B�mY%�[p��98B�)ז�-����G�1>P�f�h"�ȧ��_-���bˈ?�p^��al49T8,�����#7-6ش�=vx/���e�m���䭚���vj���+�{!��˰����)�)Wa��\z({b�_�yv
�H��$]�l��i�0���Drd��F~��&�.�����̃f�ɕ��ϟ�5d�`�J�;��?��ڴ���
={z_tt4�����gyEk�����P{a0I���]
�fV�d*]B������V}C��c8� ����y ��<��e�_�v2���w��B����]뒒��A_O���´R����
��.��W�^� �zFQQ!G//�4f�.b^u�&]5�����>��n�>A�{�D3��7�Ƹ@�/A��du����u#|p箄zrS^OG�3�5eݾE�83 �f�	"�oA3 %���#�8z&p�4�5Cj��v�$�UUU[X�)��s㭶��K�kRF�
ڃhF�����5����=��ҕ��n1�v��0���PŲ(�И�����.�������'h�M}�c3(��|R6��@v�^��:9:x��L���`�
������ν��R���X�&9LL\Aa]��'Y�JāL���������
�|�T����T����P�[P0��hIE�Y�N��<G�ʠ��̸��QQ�A��ܾ�*�jhԥ`�F�� �`o�����N������%W��cIE8w$�q���� 4�����Q%m���kD[C����������&���?�:9�t��9]-V�S���O���эI%sk����)�{i��Wިg�kHf�A|���� o%�r��9H�8"��f(�nb��s|N��aTjyv4���b�I{7���ĩ]�=���Ψ|���Ƞ��B#4S!f[�����lH5.������^����0��ٞ��M����G]jG�ۓ	�a܊�X�!�|����ݲ����4���v������JI�������5p#|�_��y���Yǃ�W����Dk�@}{��}KK�1�J�y�N�#E����Qz�ƌ�{��馶��V�Em��=_� OC�NP�7���M ��KJNEEV7|P9X��G�N�#BY��p�c��!����T�;i���v�S�pW]]]���ӯSɧ_*գ��^GK	�tJ����K�.5'��sAy�;��K\��Hb��'���^�Fxꭋ�����A�˗a�(!�f�)ih����x�Ǿ��o�Aߚ���@��G.=+쯡0���ЉM7Y>���Q��o��Aà���3��#��W��[��	'�jio7t��K$�"#���B�蠭*�A��y�tP�
ı�pC����@��<����6��@���ḥ��Ī'{w+�7"�_��O�"��A�l��^@��KӴR�j+|�"����s	��H�������w�`�ñ���'O�	��d�:��2���dQ��_�P ��J��E����QQA����Q��_i;�;�������8���0�p�22b'��*~�Fm�7�����O!ި�C��r��`���OI��
�]X�ϖ�\�?���������
O��Q��1��Gy��-|s���|�'ළ�}�?��d���Nk��4u�Ij�"�j�˪��n%Y�D�.=�]��;��������,�߅\�b��RUQ�v�À ��,�έ�*Z��J��]��c4�s��~wwi���1�܍��/�-��O��Tg�����r�f�M*U�ژX��#[�U��Wtm Y"��ȑV�1G���:��p5KԼ�}�v�g����c�z��o���O��wUB�x���=��qqqe�9z���F˱�R��Ցk��][���a�6( ��Z�Ƌ���E�a����dq�΢��Q8�ic
������p3%�`C�cN���&����y	��[�C�f��Y#B��,���+��xW�����������/q;�>:r�%υ$�-�p���hڪ�.�)���|�U�~�t�˨�ïtD�۾���s��D/����m&^*r������W�ᠳ3���,Fà3S�c�]�Q�6�K�OÚ�zU��r��"|��^N�N��J��Z��v�'GO��`�V�RC�<�|�͠��[�F��³�,HO��'�QqD���S�Rô�N��5WA�:��@�섟�c$�F�������>~k����^̐��-�G+4�_��{�I�^VV��dXGR�*��3�'���W�[�E��0K=���o������u��"�#<�P����%�$���9j���8�\�)�9@���/�p?�l���:|��2���zmz{��d��8��!�k�,+!�d�x����h�@���ts��Ç�e?�5��.JHI�N]'��]ҧ3�
��U|)��Zr%̛�ؠx�r���y�Op�g
v����-װ�j�R�E��z;;;��x�C��4��>���<>*k,�wVhn����ts�������:�#��~&;�k܊��+l��ۖ=5E����%�8d���z��o(�(#�af�O��\�#�W&n`0�˂H��'C���9�,u���Ӗ��K�76�[��nl�&̍o�!ͪ���D<�=@9%���X�c��Y�_���O
�d�{���1��%c�Nt�����s���3��]Z�0%�	�[k���ց݆BW�z
>K�/ �t;#8����g0�/��`\Hو�Ʉ���\H�d��:9�GguÓ{z{�е*8��,-�G����*�w9xm[�UZL�d�0M���XW����k/�}|�9v���wEk�줋�ǆ�[X�����M8D�~�h2f������,/..��/��Cl��XX��*u�5�u�[�������3�!D$�{�"��Ý�h8%�ړ��r��s��
k��a	�!>����5��]v��_���(SN��.H�=$����?-
,��0ӭ]����S��ٵG����h�*�8��u����"��r65%���n���U,lޘе�ʝ|ŎP�&1��V,���)�G���E��k�ЉOn��|��^<(%E%5�@�9�l ���6��bI$} V5�Y��qgF�������0d"&�n`�s��Y�x"�p�s�b��;����E���K���b>o *��W`㊮ ������%�'�z�9�O�[�����v�ݼ�vd�Xb!�ۋ)Oe�'��v׸���	�Q�>��d�iral���V�������ct��g�ȋ�}�PGl�E��MI�9��'��o*ң��x+vv{,Xʐ�a��g������X5���^,�>yD漂	� ��t��b�x�Y�5n����v��&af�E�����y��m~� ]-�ޅ����<��w�L7�Sh�3�����ĆX,P���J�T��R,w;�Oc�'���ɠ��q_� ~vn=H׫�I��酦�;4�p���R(�ER؜: ��֍��&ڟ���bF�Яu�t6�Fy� ��>�����
�VDB$��b�����B��d�+'n�P~����Ǣ�֔c��K뱛���Ő�-	�'e8$ T�����"3I�<������s+��m�ӳѺ��a��`3�TZ�F�B�R�,|'((��y�/�
� KG�����Q��!��t�7YF&t3
>����
��TCfCB��K���)����3)���Z��v�H,O�A&ka��czB:e>��c�~Ze`Z�nߧk2�Q���V��{��ʎ_�;~���-Jm�+e��%��_�hZy�aw��/L'�f��m��][�s<~c�"�A������c��Z��^�y���Z��]�v�`����2�d�F:(JKǪ+�U�-���k&cnL�sn4~^*2�<�B2wN�(Ȯ({z'��[˄�Ol���E�uY�*��ܷ��`��; �^aw�('�*2�6(J��P�{j��=Y��׶K�T	��\̨�yP��"���0�	,L�0��A6���P�n���%�k���J�'����u��p����k`�ƛ�z֭��T,���C9�� a�-��jXX�ɡu��������9?��#g������C[�������'E&�N�����|:��zn���'�`y���1.�i_1�P���G铴�ie�{����ͱ�@;x�"��`�!Nl�9�}8��~�F5N����`(_���-��Q*�n�*~��Pd��n�I�4�j���N��N4�\��u}��[`z�'�˺м��ƚ�i�SLr1�r�=e^,��8�;�*�e��M^O�x��˓���L&���e)��s�����Ċ�z����>�#���nxF����qUBk�-��[wͼ���B�݃�i�2q�W�����B�a����(�ޫ��.��w {<�󯀖9j�~��C47�㡧�CK�65@�ͣX��`wHu����n�;&2XC���߅���JDkx*LW��^��Y2�����  �b"|`��M|���V� I����m!�w�ܙж�~kN]�R���B1�ə�aW��ħ��!{*��������n�����q�"ڶd��`��7�����0P�&L��2=w�䚌`�ͬ]w}}}9�t��B��z[�Ggx�����rH���챪�[L%]��~��c�\B�a��ݤ��g�}�HUi�/_ᛛ����!pMd��&v�BvP���� Õe#�X���G��qn/���#��� �����W�9;�̽��f�S�A�&O�3�˄��DH#C��i6��򹒯�)9�Z0��K��ȒB��V+��\j�ݸu�Փ�?O��=��%h�Q'C���E�̍Aڂ�n�,C�R���-��{��Xab��v�<�/�{���#O�6�-.�D[oW��=;6:q|,�6ۛnT<��L �J���={���ңpIC7<��~ya�F��Зb'PM��g�+�U/x��﹦�(�A�aѹ�,#�p1{��R�xZ����ʮ���`pa7N&��?Lv�|�> X P�]�ש�e�l�Z�}_a��� ��!�\��\Ú�3F��.��F�v]�ip�u�!�����t��nd������q��R�S!H���3���{�����8��&�l�\qx���r)�q��DF�چ��A珮���û�K��O�;�o!ţ��$oʨ�$>���7�YR�}����
ѷ��� ٥=]B%8r ���I�,��2��رKHz!��oR��}��@>|L7�/��=��%�J���>�{��ڱ�島�.޻�
�U1q˨����6]����9U�8y����qcK�0�bǈ�,�co�{����xC(L�P`&�#�Τ���v7�y��WQ�o��/WM��jl͝gEK�N���v���pQ^m��'�K�YnȜ܎��S?�+��?�s�E/pi�$ab���Z�7�ї�<u(C&J��[s�rKmv��&�1����,�aDb��'����9g�zۮ�VI)����~�?v2��ӺR��A�V�0��Rz^�nfk��J�$~E��/d�ކ_;���,Zs�k�l�<ޮ<�V `�B�kW���l�&k��Q71���{��u�jۈL}Ux�Wr���X����T2mJ���4T�Ԕ/���z��B��U�3/g/�kV���`<�g�� {��Sj1�Q��%罔Ґ!scX�W+����<���F4�R��RR�����{~{��|�~~���>��є��E�!��C�j�x퐏/ݤ�������Lf��L���m���X���Y2��E;;�o�ꬃ"��ܾ7V��ڟ��م�4�D�ѐ}���S*	dF�P�q ,��$��ŋ3���c��Y5�-R=�Xl�����V�o]���+�l�]�B�5<�e�Q4�
�f��[	KX.�/
���eI�B���(���P�'�"+��.B" T�bz��^rE�e`��=CDU�h�0ǃ�F���aU�*c��At�7�ևi�b�-!U�w��Xg�i_xd��T����{���,�/H�Q�ɠ[�Փ�z��Y�E��a"p���W�An������?���c�E-�.6�B>��I�pE��VV��@�=8�P���)� ��kY�
�@�rz9֛���B�$�Uf'K���T	��"J�ޥ����}�O!�� ;�b8�
�*�m�A��M�#!��Ȳu���T��+;��e�@������_ L��µ�Bڦu�T�R����s�� /�r͡�N��6Q='�u~XQ�����
+�&�j�B�4�?��Ȁ	1"�(9�PA�T�!��ν��4ϱ/�h�:��ѹ?��c�o�����E{!������-v��Li��MW��rB�0��u�>(���.h{#]�K�+����;�wuD`����E}2sEk� �,��ߚ�گg�"� 3����]&X�T��G�#3�N�Q&�E&úU��@�����E@g���#�Q�/���N�)�����K�ݯ6zd���8��uT�(2l�ձ�ETok��(Ah��x8����Tg�|Bi�@�܃���RRj%�F��l
�LI����-*�����S����׼hR2:�p����\B��
})�-Q5�	-v{������D�jb1�x��@�j�U�$ZD�kAFYꉄ?}������i�R�m�SG
$���_�m�F�L��2f㱵�k�s?o9��M�"O����,DkM�կ͞��P����&�*cn._���<G��\��c�<�E�<!�I�nIMM��D0�<���Q�h�/7g/���Y�+̣��A8�������� ��0(�z0h��%��s���;��ɒaø�{l�C���=N#:���d���'��̴Q`�Ɣ�@LI˜�Vf<Y�-I}�S+A�Vgy�'��*8rc�Ҹ��}(�^�-ND^pشdk���Κo�?X��{e�]�v��]��s�[��7 ��s�a:��Km�3��D��M��g��G���eB>�a��n��<4�;�4û'����N�Ů0�#��b$�R��c:��zU}���6����]&��{�����Q�g�*�G��t.ݒ�_@�Cz9�TjFR(`��y��@�Co� ��y�q[r�0W�٤��E(� ��Bor-O��@OG`p?\*�͗��t��ڄ�����^K0�-~u~�&@b݃����H����0m#ݥ# ��Ijcd���vy��Nl�XS�~ '�vF:
��Nё)�
M":�u�[7�x{#��ח��d{(5"�;j�uCk��j�A,F5�DÖ!8�uk/���]y�))�"����XE��))S.�IX(��'S�ڸs���9���8��$��b.p_���71�o�ޢ]%ɔ�/g9�q㑰���t��F�}݈��j��	{7����<�=��6�vԙ�a/�W4��9�,p6;F��,�NY�L��C�H"�10�gv��Ú�yO49��8���W ��A�1A(( NOBuP�����1����?��1�v#Je�<��GO�B��i :����sB'�2|⍫����GE{)	���$�8�}(p��%�#Sc�
(r�ؽ�#w�E���4Me��
�Η�A�2����mB��!l�aaЂ ���,���3�9<��:��C_�f���`7�\2�RRp��O���޽Ϟ�>�Mݣ4��� "\O�B�9pO�k���^3��.B���M��$=�u,��hc��I���K�J]J��:� �މ�Ԏ�[�J�ch�H:lV������}[ی�v���A���0�ފ�X�� SJ�	�_�2SR
xM�A©�f�	�j��=�Qs�4��E�0~g�&��՜�;9g�L��EŚa��;�Y2cA� vږ���k���,��:c-�*T��^,�0�"���ee�+6G��s�5'�k,�x6�f-R�&/x����~�s�>� 5q�����@��X��Kg�B�U2�5r��۳̀�t ������ބ6�̧���@v�9��-4^,h�����Z�E���uFL�Jh�C�7%C�L �P�!��f��6D�B�@���|�w��*u��olđw��uM���9��"Jr���[s@��A��f�u�ģ햋X����7/L��#��t���PJ#-������Pv#���h��b�M.�T���If����9΀�KU"��<R�5�2_����W���P���U��$���e��A�i���~�ͬ���	�̿At�g�vE��sT7��0�J2�g@���}6B�P{{�:%����х� ���Ċg[�%��(̾�rU�"op%+��-Q��n��* ��틸R��1!�ъe���u�5�]�$daiQJ�T9o�嶍#7��3fDjf.�����P��)��x�&G˪�����	UHf��[�ѭ�X*/��)��U�"/
�1��t�zz
j����<1)��lX��"�}_���}8Fz�h�S{>Ta�����fe}�@�O#Q[��ezή5ǜ�n�[�B]�P�2��|��xb�r����/�M�TP���Ix�m>�����j��<�-�2К*�"��J�וރBp��9'û���U�����s֯S���'>vY.�S��U-�K�F�����Pl֧6^�~Nv&��@���*� �G%��{y�>A+���i DT�F�����Ŋ�s�Bch��.6E�1�l��{�ӧH����&��:��B�e��9T��í�|�ڨ�0�$i��:l�k�Y�o#J����Ek�����b�B��:����_�]h�X�y����@�g�Ȃ���ݪHSl���r�e B��nrx�4�-�3H�B��]��HI��慺6/��+e��łJ����2�f"��@�+�T�����N�-����v���O �:��-��}�j�3�������AJ���	�h��$^O�h!)��>#� y��+�Q=�ѧ"(q=�[��k2{��	�Їӭ[��n�ГAbx�	b8 �d_,9>8\s��ğ+�px8<]�^p�93�!�W`>P�򂦎Z���\�(�l׿ї�T#voDy>s A�Q���,�t����h�a��&P�E99�|6
Xb�����XI���ahF����@� �5��.u�FyU�$��jbà�7�$.�{Np|��LFX�ٶ�|�B��V��A�G����wxRJ�X���GM"�����r�r�?6�bM��tI")\��޽��ӈ�h1��R�T Ha��ޘ3�͍t�DK��ܱŔ���R��H�G��[2��<����yM��m�6�[z�B�߀-���#���W�h^�o&��}Ȏ,������q;.f��q�� ��RR����޸�R��PIU�Rk�YpǸ*��.�����7f�1c�h�}����	1P�11_QfWd�Z	P\����m���N���q��Ե�ի���ߖ1ӝ�擲�D�KG	��@J�[(�<�J�Ғ#�8��/�Z�f�@g*�j���`��S�iG�q���z�������s��j_1��:�CS%���ja���T|u<8\@ɼ�a�y?��M�%DG��L�_������N��Z"�&_��'L~��F�H|ˢ2�xwi[�W��p�_(���aY���w��Q&��ZT'�{[������Q(j���k�������L'�b�h�ƴ�4�ˍc�4[Z��#ɘ�����4�m�S�2G{��%��d�����"Cs��ڇ#8}z���LeJ�^�'iR	<�`xz��ׇ��mff|9T	s��k��D�7�f����ʶd�4<}�H��baK��\ZJ߈vK�.D�<.�Tnh ���3+�{v*E�%"�f箯��r��U�!(~�����":�()����9;�>Fr?߼0�8n��+��{�Q������� �[K$�ؐ�oAD��]�F�	�횃Tx��X`|�6R��'����4��bv��4 ��O����z~j�ō�A�U7̝D���ǿ�datLdr�G��k����)@0\#9���$z���ȉ����KԀ�/P)4� �K�K�d�����w�y������*ꤦ|�D3KJIф\SD7���-���I�d[O�PAUu�Fy΃-,$���1t�[�r���XE���Đ3�m+)�ǐ�\�C�^����@%��d���(�aX8��Y���yDKa�y1�⿹B�&�b��W����A���G!�� Q��B��L�Њ��#g�=�u���ۈ�3K(cÏa�d�g��$�	�;*�\F�LV�:0rj�O/O��Ff�w���&��U1/H.��qr���Nl뱡{��q�oJ��i(�@�J�|⍠����O41��v�f��e <�P�n�I��pBV�D�#j
Zxb�W��@U�B)J�fba0�XJJ�o'^�DB@��P@�̡���������?��ڼ�ī�H��}iD--BH�kt�5�x�K6�T�n8��r��F��F��3�-J�) `���ū���c�"M�j�Ry0�8hi)"pE@��!{k���/C�ՠH z�ӆ��Ow��5�g��l��Ql���1�)y4o�_`��|�B)���;�Ġ��Ea%~���0Ū\�:=E|'�'��P־|>h0<b�t!n��<��n��%��k�~�
۩m��aK�����ܡ��	"��������b�w����k �O��JZ=���-�Q�3,x����\fU��R��%�]�-��ù|�Ы�gx��e]G��aySD
�Z�>�yM���P����}�d�úsPH*"��&O��z�l͓���+Nq�{�\1��)'��_L��=�ɞ}�����V��Ő퟿"���T�SY� R��Bp�a�}��	��AaXR�Z��y{���"���c�D9`��N������tþg�#f��o��RgO-�1�NhLkN���6r> N��qWP�����X��b�����XX�^[�Q:�B:bhI�҄�t�(��#��w�?@\M�nr7���>v�!T�A>�.�k��m�4{^,�c�� �?�AJ	�����BZ ��dJ��&p�W����R�c���6�2?�H �H�)
��
���jQ��XzF����M���V��c�T	��(�P��S1/��+���V�S,�(A�{*�p���Dk�EQ�?B�C�,D��GLiV��^�i��A6�ҡ<A9er�J;1��j#��E�Ƃ�.���!�颦2���3�[|�d��=5��{�Q>�����n[S�^��tA��^�!,f7J�����K�W݀N���X`���Zrü<6[c(h����Dx��(X��%J���&��f�5�l5'rf]����it�i���!��1=T��]ʓ��QL��.���rSj��]�Ҏ�Rw��J�Ȃt���s�ʮU��s^�J�ɡ�����k�x�)�J|��Mtf;��b�E�ޙG9|a��Hp9��̮4=%r^�5g^M�K�$L�	���ל[�����\��%:� -.��%z
������e#d��E�����܌r�5-:@�7�Μ�G�&~�76��R�0�Yy`�M]����\)WVn�]�<��_t�~}�.�j���̶�α����U6I\t�ٰ�@4�/2�Kп�Rb�Z�7F�7lw�8k�3����z�����~�9_;����,�w^ ��m._��I�P"p(���3v}����{��p1{Hمr�RB�7a�'U�y�乙d1�g����M�ްz�w����hhTR�2Q�=��w�J�M���1=;���Gل��T�R�JN,�h9����I���va�6�'�#�؄�~��k2��ƶi+�	a��J�h�f��Ϝy'���5�XC�X���2�f}?�N�k�F�ܓ�_I��N����u$(���ޙ���m�w?i���1�I�Y�
�R�[C��0��ӓ-����~q�����fʦ�Q�����,�;*�/�h�{>�����a��KB�oUa��9���:�O��f�3�_<Du�������ϸ��|�U�k��$�;%�z�~
�)ﲦ�m�f�="/$�\;�y��>x[��5i��b�x#�҈mG�{�'� Q��}Q��DW0}�~NiQ[����oJ�s�)�?ij�A<���%��B����.Vi%��Rz�Vq+nr�9�s2ւ���M�
?�0� ��<je݌�$���0S��ɏ�D�����<B��-Mw~���O��]�J�_�F~�_��[���[��[�i.\�W��w��m�.XDQ�q�[y�H�j2 ̛����Ckm���X�b�:��I}iz���Cfˤe;A��or�c�f��[]uߵ�L��g��V�~�]�f��=>J�̇���W�g��j![,��%a��o�����뉕t���Vr)=���1�1<ہ���V�AF�;W�u�'ӹ�@��:p�*��4��;���ۤ�9�T��,����g�Q�{h�!��ε�;L��6r�
N>Q�~"x�r+����H"JYb�Ȥ��"�������hh�ۄ���-Ӭ.^X��7I�d}߲L8��8���������)p�9>=[��.d��UEe2/��������?S��f�m��0�zb�t�~�����؅^��Hp[�9�����\���T٭D�IѾ�%��ғH�4U��]��E�$��$�$�r��땢ͳi�<�\&˰%���V�%��.�;�%��z�D�(͸ub�7��J��O��ʡ�>
�����z��n"���F�OYm���qZ�Ή5�-�άƄ�X�k#��ȘQ��5\"D~��:�}�XJv�d4c2�&�ˈ���W�d�*¸?C�������7����`Qݜ�$�;�Efx�6,ʝ�$�o��b	�#���]Xk����S�"?c#d�~����E��lլM�p�O�ƣwF'l�tRQO���B���½�w�p�!�u�c�O1�a�CG����Y�ad-`��գ��DV��"���D8*�(5��5����b`�f_�[x�N譄ӎ@ �W���/kV�m's�f�b�0�9&�-������#)�S25��I����\�.U|jIg�����s(S�����\�b�P�	��i8�z�^��T���{��2�M��\\/�0��h�Á^�e�w~��r��4[j��=�8�Heb�ף3�	�G�,�Z����6�,)H�N*��3����?[+�"R<^I��d �(����*�����:��b#`8��⩋B��a�p��)��h�Pb(���D ��؀�Cirb�Q��g�=�2D=rt��k���#���h�Ϣ(����a���ZVc^�lO��Y^@�D\_�����?��̦d����2,V}`^������tl��JG_},8������l�p�A�Z����Tw���I��`˻�)���֬N8��5�L|�k` ������#�qwҲ���2LC��ېc��X�	�C���74���^��<A�Epwܖ��� -��J�5g7,^��I_Dq�X,���'��*�S�>(YX#�!��˧���'�7T`@���ԍ1���!�K��*ޤ9Pg7k9��I�h"O��  >Xߪ�d��ѝ�E{��t�oM���=����͘'5����	�*P�:ݠ*�Ҿ+Ӿ������у>���42����X6#[r�=��܉��zS���/醢�PP���砲�i=m�T ���^��y���f�_(�}�I���
�ӫC&���_�1G���w�7D���Q( 2�^��� 'Ǒ��"��-b�M_b-��'>0��h{��e���&��w��#�n�6�<Z������UNa�t�ee��}Q�T}�̽����/w[�gK�R:�R:��6�q����D�����]�8d.�Ec��R�葄C���μ�
IN/�`�9<��`Mw��w��"����M�*'�
��8�m��?�l�#��Y�N����	isB��4�g?s�vH�)� ���Mɇ��w.�����s�H��-I���PZ���q�<�N��K�͠}@o��v��)�"�KϪ$� ��[HeS��b弦����=s�7
��Џ��ӲeC����>y����2��TQt�Џ����x�DVq�V���&������1mM�yх�7uIs�^pb�6%�.�w��b�_���5��ˇ���ks�c��0<�`�������zJ�K�P_���ғV֣ϖ
ΜE�_���#1�]��V��hY�װrm����������d�;i�*�̠ٜ�Z���FSk�o�Y�,�E��i�P�saY�3)��#�5�#^����p�]v�G�x��@X�+z,�E�b8ڽ����k�U�u��L=>�����M�@|�S1{�'��K�>�PZc�_o�����0�w=�����#*}g�� !z�[����m�洠�E� �C���"�i��C)�м[m��כ�V��E�
�)��a�䂇�	1��?δ31o��cV�W��t��>7=�˩Aˉ�Ik,�I��{�I=L6���	q4@[:�>��&�ݦ$w�#S\u`���L^���^`VG���i�E�{=���ށgk�(��n��_9R�Y|ta�K3b�(��2-Z��\����#V��"�����2����RP�d�	�ю��b�W��:7�cRЌ�AF��V�[�C:�?��@W�#�U��s<�'���_vOJa�W�z�����R-�w;U�|�R����
����+�2���	��
�t�c.?&R���*"e�u����E=G�(ׅ���Y�����P͎�&�T'9w��awH"9�����J�ag���1)��`=��b���`��Mj���j�䏢7�c�{TF�t�ؕ*���+81!ăH4�|�%S/��������g���`�M�c1t����=1�Z]�J�m�E��ߤW��`�0>t�&T�d��Af�&Ν���]��a���q=��7Zf�d�AN�t���B�o�:��?�X�D%�%��:����S���g�,�X����#w'�Vj�1-IL$��6A��������� j�&ws��9���W�3f[���T�:��0Q~)@~�͡o�Q�>�E>��|�7��yơ��(�؞k\?q�G��
4n+�B��`�u�"~k��2��=�f�����?~:W�׏�Q�h���%�a08�����.�W�ὶ��7k��>+�t�����X��}��O%��2�r�I7~�N�O����n� ;}��l�S���k����s%��9zT�2�<m?��!)�u�������wI뮂��ڴ1m���}R��г�-F�"^S咨�Q �X�� 
�(@�-�����Ǣ��f�i��齄�d[1��庣ia{�FX�����=k$�pjf����A�a$�0|��""�B (Ķ����Q��,�Pb�?2��)���-���tP�^��&��<8���]��A��5Uts���tG�L��v{"4��{».�����׿�`Q��U0ڿ��-��}·5ҷ�J�Yq%,��`�G��cR�7�8�L�u�b��=<w��?������y7�}��Ӳ�,,���Do\jf�fj������L���7(�u�!��.l�ݚq��2��XƳ�d�8�{v�H\3��O��n�%�9�%\	�ɪ+�L�C����m&������E@��*uT�FS���p�2�x�)��$aV��]2OZ�k��Do��e^�#� ���=�a�0�x�=l�JZ��т7z|�C�sCF���L�/Y(ȫ��wܜ�]\�����/��K�"�m} ���4����?��ݒ�iYJZv[/uX�4��q�d���)�C��W֗m'��!�60f���y���,�9�u�x���P"썰L�s<v�-~���W]�{�Qt\��{� ��W��}+���6��Yf�%oN��C�8�	�id}ѩ�|��Mq����~��R�� _���1�O��"� F�lP>��P�K���UH����4�{V\�%�2�/[;凵��_Hާ�}���W�^<�G�����iO\3�:�i֓*_�hį*�y!gxs�2��iECa�GC��8�������y��Ө����~���S�%F����ע�zCsZ��l�[.J��K
���7�e�.A9X>`��1߃=$_�(/_�jݐ�鈱��2��.J��_�����x�����{S7ѽ����ݨ&K��n]*��U#�ܡT�d}ZdK�Ie)B2b�F���${��[��{�3K�������}�ky����9����u��R1�Y�ʪ�.��$:���}f"�,TƗ۬��#�9-?X�ً�o���S�ş���q&���t���P�{W>]x�25�����Oz��AYP(:N���h/x�$z` ���q�� <��??��� ��h�|Q�XV�I%���)?�(V��	�_��\�ĬF��g���aF&9�|n�������0n�~L8n�(�sUvu���P d����4�B�8MQ���v�v\�ol���[�;��D=�s�`���\܏Tt@����}	��,�|g���2F��q!�����'>L���v����TV�3�ƶCd��C����?�3D��%k�Ь�2-��;Pg��u��H�1�Ч��eʔ�U�언�1�m2,���pzɇµq������:�8������߼�i�A�[�"��Ҫ�f�	S�f�q$�+��xm���g*�z��v{o��n��|�_^=��;%,��(�J�A-��7,����)Ѵ���V�zAƈ�����X�U4���a�{�[���ŝ�l���h�%HA'Lx��M���p��%#���8ytY v�ջ����_�C'���c;�<h����vo��,���ogw�J�ݵ�s9�aK�%�����:>=�:���-�����Pʏ>qU�;���v�H�7�����r�[T+�e����0
����.�w��\�P���{]h {�wj�R�+b���8��^?xP/�������\�	�Z��oމG@H�N>g�yn+?e�6���IGcQ������ߏ~��b�8ˇx��(a�2�쁫x��n/�����~�7���g��������;�xIc&�(�j��5�عk�Լ[�e"l��3J-2�L��1�TlDT���@���&s�k�;�jZ�'�ۖo�#�$��#�AU���-��fN�tɔ�Gզz'!Q�����|��E�<2���]F�O�nq�4G�z,?����Q�)��C�;+2�=�]�����_4On#|¶rHn�s��<�S	��Tns��<��/�����e*�S*얃StK0o՚��M�y����v'�a�:��:Z��j�Ӈ2߾v^��2�1�4��?;�>�8�B+ϟ{F��	>�6�dՄ�����0!��~�[�H���6k[T���>Rg����?���fi�� ��a�Y�s;�~s{��Դ���/読���I+�������\W>R��.��6җ6�o�����t���hU-�����'ET֨�%^js��{3[�]�r����G!L�$�J7���fq����
o��������2�[Y�r��5|��~���'ܡk�@g/�Q�^��)�K�!�v��mxT��d#F/��a>�������ˠ{�!� l�r�@�IEFF"���K��/>�\�?�Af{�31
V�UQڣ�y���x�8�[
��q ���?����n�H��Y͟ϧ%0逾���1��X��8�!��rC*	~K�_�t��
�'�����\��g�&A[�@�ۇ>���`�F����]��k��`����֋h����!U/&8m�^�88Nw�p�=g)��EĞ䎛��1��{ǟ�=Ϩ��Ƕi ͡=���v�-�9�Y� _�:iL�Αr������f�8[Qt�G�
BԢG(�ooq�(�4�T��w���ř�JrV��页N��{��z%�6_cCuh� v��N�h�5������� ~T9(���ufF@0/*����F
�t��Cg��u/��Ƅ^�i+��]��̞�����w5g�����q{���n �_V�`���}���/{�C���K��j~'~�P�^�`p�	����}�J��x��hi1A���3~M��5�?j��8A�Q:������О#����3ɝw���*����e4�{����|YK�xf���ȂA�}��5Z�1�x�V�{�x�ۇv��E67�-�%����:[3���
j�_#37˖��e�A�^љc��+|���绅�7v%�Y)�H�]$��V\Y��;���"Έ�g��s�����.ϖ��*�f��:W�3tz�a3V�b��
[}'�7��~5��S��+��w�Q�z��L�Õ�:H��i���?���v||��l��v����3�W_�z&����+�܋����P�D(��Y6��1`O6�w݀�1rɺ�Z��33�=�M���WN� �Aɯ�w��{�r�$�n;�d�J �����\�Aܿ��n�7JH��jqlɯ��ۆ� x�qr�3�����4��,����Ƀ�3D�V�]626>~�g�n�oӳ����W0m��6��ݼvp���qr��[��ttt�<�Q(���5�y����8����3բ\KG�[�7�����{K�y?K^4�w�.J�r��vWa�%^�٭g�Nsw�q+����0�?{�`y���Q��MSS37�_��VC�d��Y6ZXZ^ o :v�hR��rf���������`�#��K��p]H�Dg
�:	0�g�~@O�o߮����F�p|LR�q++�����y�h)4�/���7�󍊈�TV�I��T)K���mE��K\Nh�G�`544��/	|�?F˟\�����<�
cŅ��w��޷�m��8,�:�TW���a�`�B�~󒕕7o���<�������^^l�nS�C^���o۶@E��}���	��U#��y�ɷo��z�*�T��ed��)����SYw!�A*���@*8�^8/wYp���}}g�A�&�']�2�!L�"��1�C���ʏG�C�y�ոp 8��}x��?�g�� �RR�{)z&jaGɖ� �l��߄��%��,�)��I��W��&�xOu��9X)ӌ?�zwo�9����oPZ�=�o����
W�kRbl8�~t�¨�1�>������k��;�	B�"��ޒuGS6_�)J��g�4F���8!2**%��7��0j��#4,l�^-�/χ�� %F���W�<Gg�j &�2(^�_��R-7DY�~�����ᖰ.���h<D;��U!l�0���q"��~��\��8��Q¨
��c���22^ەm�������c�-j�aP��nn��E-���p$�0�wPY%nL'�	��vZAf=��+%�}�OM���7��-��;x��Q����e~o���B�@XVm5�H��ZX 儷�zSB��x�!*�Ke �Ƿ)(�E�v��M�ܯЪRüL���r����8�{/hT�h9��'<�PSS�0� �Z����7�4l o����%^�G/Wb��74A:��^�y+-%u֎�S��;f�?��+GF��	����N�M�aPP��nѳ�C�po��R}�֘�ty�ѝ�B�ah�L����5R*~9�V}J��hSj?��kU��P�}aM� �DT{5mS�Ȧ_��+E$Mm��!Jlt��N�H!|�������w�⇄��)�� F�'�OP��i~���+G:::�jy���NKo���ĖE�f��`�_�V�+l�w�@��w?_o�GRP@����`�E�{�:�15~H���K��|��xzf#����'��֏�w�F�̈�LTd�9��AQ-Rm�kC�;��b�|�w;��Խh����,��M�E~���ٳ�P`��gS�~IY-bE*���.��Il���uhn�8W�cP&�lݺ��J��ᳳ����{��,--=	e�:�tqPP��c!EWl��o޼��f�A0���Ǧ1r�R�L��&�������?S�G��5�O� X��III�m��7Ç��9�}�`�S�������G��F����36ZW�\�����ڥNa0T�Er<���K^ꤲ�x:�k�[�q?G8���PQ@Dq�8#7w�xT�$?�mVAT�8�E@T�����C��^�z���mTW�`�!bbb(���AHnÿ�A]q=4tP��U�tt�6��dI�Pₕ�Xq��u�c�LR�Keu�<��Hz���=��H�MBB��:��?&��Y8�aF$�V���ݻ�#���75uu�4�/��j�݆e��V�ɯ]��!A�9���W�� xm��~XI
�J�8�� l��^�Qȉ��[=������Nԯ�N��:�E]�h�����Ne�^	�f�?v.٤��o������&�w�6��wM���;�ĨYH���� �c��V�bT�`����	�O�IYs��v
Ӫ*./Gإ��p�֬��3=�/�~�/xxd��}��@@��"�1�i�U�����6��#�;65��3�Z8�kC�C��H�̤�9*p�~�7!׹�X���3��;9$Ե�g!�B~�RL\<��8�Lޜ��Vܯ��oq�M Pn�|+� ��1�o-�J��/j�r��v��A'� �)P,�Z���QN�-=��
(�K�@�v���6�_��|8�����0�.��z�O�����z9y���D �08~j�?BN��eee�)�I{!!��P�c�6_p$=jw�zwJe� ۉ�UV�$$nhۃ0���
4p�d��&���1���y�%��)����$��V��0)(ꔛ"� ���0����y��ֱ;w��C�W1������]��!�\B�?�DK�cP_�q8JF��0��&<�(s�A	H�����qU��2<{��'%%%�C�_�2�5�΃���Nw��f��]��Cm/�[�(��7���9�ԴV�|��^؈b'J<B �nX@�hn>^߸��A�����4�h�O�}=:�ޕ�O�qm��O���=b7������u�ʃ�B�O���_�X�*���oGFΓ��v��(P�QYU�?8����l�j�%��u!�7��x�-�G��B��נ���~����Є�/a��j�yf&�zoG�.%��6�Z�2�[E&i5ȹA�C���e�q�"��t�]��\~����PW�'#�?
�h�F��+M����=��B���0�L-`m�av>`�p�������^kQH���$�777\j�;�����88�Z4�K"��D�Q�����jh������+�H����;��	tĀ�Jf��k֤�:�w���³�S*Q���B�=x����I����޵��TeX��_DDD|�"��	"(�6k�k�[9��9�1�>=��kzzZ��1��Z�I��O�I?x�g?>'~����I�T�L:�i�-��x �s���>��m�"�4���yV	�P�u��8��1rLt��U.xY_��}:"�N��]�Gq��~�<66V7T?�6?����h�Z�@�;�cǶ���,Nh���`��	
���W;�;�f3�>�����5�-b�#��+�Fb���¥��Qul�I�C�RS,-,�n~[�8�ڝ�6`��|owE^�(qd��y1(z=	�P��[����]�%�}PQ���/�J�px�&�Cx<FNJO���e/�|9(SB,����g]g�D �6��aq0r85� Mb��e����t�;d��}�y4f#^������C��%������]�=�3 �ǈP���t�@���եIe�!��a;3oUH�u�j�,x���tq�sL��:v�^��+;�I�j�Jص]�[ߛ�!]X�{���?d�l �==bY������Z��^T��Di7~�X̫{$��AG:+I��P� z��Q���p\��ʊ���
���#4^[�pwH���e��8���O�M���������]:N��{�.9�i�D��ދ^�qT�$~��Uww�8�S�(������f��P{�vv�FG,��A���������rx�}"�,��-@X����1P��޵,��E��__��9�D��r�aEu�c���GL�ʬ���I�A
Vy��9�x�}��ʪ%�t�?�B�MM���kl	>�� �pB��~�Y��8~i7�&m�����6�jj������Ux��9кT��E�����Y�?qb<\Z6W6��_'�%�իW/W����l�����-�L���n�@uxF�[��:i���q�C_�cVfݥxF	"��S��੿v����v��jDQ໫���÷�Z�lװu?I�@��[�'��K��D�|n�6�������|�<+1W�l���f8�Z�����靐�������W�z7s���b��\[绺�*P��P�7*���G�� ,�R~�sN�[5S�7М�:�ln��)��\�0�9����N�u-�n�O�Ksv�����D�qο��
��{���^�뽆��[�q!��f�5%)1	=%��y��D�Wj!��w�X��;���@}V���z�l����7\8`Y}���Ԣ&�JN���(�~�kg*9m�3	[�*��� 	u%m��dɒ�z�J,L�����
����qc�[�j)z�h6AUE3��M�n�����X�s��L�8Y>��o��t��j���Eu;�%'�-��0����P��$���2���m7Lq���ʭ��l�������f��6����㭾�p�v���+~��%���0��y555�q�(�g�:m �� ==};[-@��7�?O�B���҆��Ĝ��(�1[��0��^������a�oS] y�H�u!�;{����$N��*����������\�mo�p�_7:�H[4���g�� ��;)��ٝ��_G`��R�'I�E��F>}vj?�Iu���w�:J*��zA\3P ���PW�OH�.�ѿ˥�N�]\\:?~�X"�d���c�����}�qF\�f�h����4�t�A8�رc�5�Ø�\�0��}էTƧ�z�I�?��F&2"��6H�$�����2Fߐ�kf����η��s�ţ~o�R�i "e����>#-�䟆��JS������v�����;�x��̟粆��n���pY9�t��!�5%��Ep��`f����<,��p��k��<t���'�$1�^ `b=��NB>f$�w����]ZU�|�7����W���/_�n�˃l ���\�j���2,�B�t��*J�r�9?2���i^YQp�<�m]Jõ+���e.�4Q�/>� �--IP|hj���a�Ď�=j���`U)1ᓒ7�
�>�ef��OM%@��_�P�]x�I�K!GA��c�ⅾ�=��.x����N ��1r���6effƟl��Lf�LLC&sm��F�(}r�3*+��(�L�ε}��U a�R9��ӫ���S�	�!�0��q�w3�y��ap��N�]�-���l?X߸g�:��t58�e����99ڥ��9p�W�S@�Y�a5�FO�������7�d���\\����r�P���!�g!����f!ձ��\�S"��~�Hs��y��o[��)���r�j�T�*voh�@���x�8T��ǧ����ʈA��c���!Kh�_*d  ��RW�y�k��1�q�G@6��X>�y,iKb�X�K�}F^�q�������혶$��G�kO����T*8̗Q�@�+h�ސHS-�KJ�:�3:��*L�;�a�,D n���������>Y��<Hv�f�Q�$���-k�?�٢W��R��Ė�u��VKl�O��ȼ�����߱�������o�[4C[-�.3��q	q}%4�֎�J+<x�Fӆ�#�q����a�{��FG�z��V��w]Y�gO��&���d��F*�*�F`*����C� _VWW������y-Z��}��3^�<�,�o�Q<���m��:�<[��?6U�H��F1��(��(g>���M�?�a1�'����;gTV�Fك�k:�u����i*���ഛ�cZ�yLG�/$�����"(���D�h#+����|KX�JkP���Q��§_�f>�/���r�$�w=��Tú<=f&�� ��"�#e���b�2�7���9`�Z��N#8}5�_/�+Q� ��*]��(��R珧���EA� b-s3�Hd5��:K�25ZUHh"�m\n\87�[(��O��@#��'+-#c�2J�*����4��&��h��w;�J�6ۅ[�����8�bE?��^bo?�,V__�B��r`b�H|��
Ѧy
�.�r�v�_��	盔�Ѯ]�gΝK�뵨j��!7�����j�Rn�ٜ�����	�m'b��v�
$��
�*a���~�=�s��?pE`�d�ܝa��)����@�,)_�nB�YW�)����^)j�����Bא;ɽ�k���	T�`�;�cMN�|��d?�������~7���������h^�Gg\��{y_���E�9p`/��_3��H���|�ʕ��beϋ[�[�j6��4�$����i��ܜ땔�< ͌���~����[|�׎����@�;��̞�k��[�"�!I�727;��� �瘸d
�`Д��4S�KYf+5�r	J7~���FR������s�)'��p�KIK_��3M�=/�>�:�G� �9��tT�҅ǵ�VΌp���&��(�;�zo�K����| (V_�:e�e���P����<���=˰H~�;fʛ"ףt}��L$��>j� 榬�T��C>�X�.?C!_����p��=ē� �AP�����]��u��[�=(��^�^����I��U�i0}C{{��Į?ny����r��6p�7ڲEX���G�F�燗�f�Q-`+Uz&V+�A�@��_Ҫ�WǗ�F �&�'�J<�ZΕ����')Za��Q�PtǛ۲z�{o)d�4E(gtJ�v��l��A�����z��Ӡ�'�����A���1����*��7���;�� ��=��\y_O0�f(M)����Ȑh=��ɀ�xd�
�/�mz�RƧgAX�3@���7�o��+����Y50$T��̒[%sss}���z�k�����"$WB�h���C�?�*��L��m���-9�X���5���g�ŋė67�C{ZB�@];w�1�z��&���|3�6�';;{�]| \ �+@�"�<<6H�+ǃ<s�L��De6X�_?vx�c0�crM�e��Hޱ�[$�LfЫ��U1y��q�<�xx��P�?�%�p��{��PZ�M�"�-�@r���"H/�V�?!�N9<�ַ2�hR�лɟ��Ȩ(sc#���e�,,,��hy�Ѧ?���>�6��;p��7o���/ �Q1��Y�4�Q�^vMsB �|�����V���>�2�|9ȟ��Y.�h{O<�D{$�����=c�Љ&�����b�DM]}�,]�u�w�VUqM�qP��m_�E���W�>\�0�݉�E0�w��{�#��?w��f�R�V�t�������{��jOgX��'j�-������E��Ӊ�mFo+*�V�^M�������1^ T�WP��cp��I}�	5�x������V�Nl\�3j���Iڪ�a S������#Y�%WN?ѐ�V��+����xL��xqw�i��Ҷ����̳��W쫢�icp	S.p�BS�Un��R�|+�U������;jN��s��bP��O}ێ����Y2����ADՂ�o��W�}Ǧ�u�x���Y��>}��X�x�u�_/>�'��m��:E�^���ϟ7�.l����l��]���6��R�Yû��m���۳�6ˀ���E���V���eVN<�W�z���j::b�]��O����6��X�~TW{�`�VSw�[����\�/D��(ơ������V���0K(����辩�a0�#?�Z8?zܯ��u�Pj�q9ާpv'�,�P+T�H�;}��sSS4���#('��^�}��2[�H.�*�999���uo�925ȦبbQh��g&i�u���c��t�P�rZ�{ �
QZm�i���ҥK�Rbf�0jB�������I�@!��B���� �,�6y�&���C�ìƥ@b�S������Q�m�m��se�TN˹�[�J^�zS $����)<ɂ��Z��OL�@��"�v��(\���x�W����LQ//�Gr�����G��[}�#u{�����	%���0��+eV�VMC���D�6#mϑ�8t7�3(��5������@Ͼ��т���55���ۣ���uXJ��U@D֩���{��ϗ��e���t+o��yP�}d���A�����s�%^��'����|�ِ�U��sڮO?,��D/�}l�Zi�o��]�%W/�8��H����~�y��g�"��4[�+�|r�-TM%Mc6��R�TCV<�c��o_w��[��(���t�p�hb+�III�_^}���C#�M����Є�Y�K�#��W�� N�~�yh�<М�ڋZ>y���l �A�� �RA"<�]-�|l���D����&9Sw�\�]�`���d�V�P����щJk�n&�Df���Hw~y��}�V���h�A܈,�T��}�b&�Ҷm>]�&iŊ�9�%)��O�A�t|�*��to4���j����L9��b�6{dnL�ʖJX�z�Q�r�(���B�)���c��Z�ص旾�g�A������uuu��ㆆ�%��wns_�xHBO�>�V��P}pTFFFj��t6�h��������T�ng��r�6/|	�2��?��OYUW��t�3{%�f]�3����o;X�y�����#��b
��-��,�i7�w�!�FÇ����ǟ���"�������r�6@?�W(�p�eS�g��_��f��E�l�=ץ����k�Ww>9���y#Vc��q��J?%�U��8�f%(�������) ��w��Ѵ�W][
u�F�uf�2��g�����ɝ�Y�X٪Q��k'�U��Fe���N�-�B�dl�Z砤�饯ǝ}+��]�7;ɣ��Hfh�J��#Ҷ���a ���|�����o߾����~�#}�X�h�o���I�t.���8�Ѵ�+�	�+���rfpwwwօ��yks��v���j]h)Ե^0x	
�;�u�툐�硧�1���SI����PZ>=ޚ�刎��[�����J$H�����LU��T�m��I,	

RRW��b�"q�=zM��j�7z:j�K:�B�]�EG+�Zf����wF��ɕժԈ�zy�������߹{�=|�LJ��蘻U��w��~���K�j�� ĞL���MUe���ٻ�VA��z�*���9`���k�R�D.�ٌU ��Ρn� ATa�~KOOϕ<����%�\�\����*J;�(�6<�bf�۳�<l�k�gt&ill-�=�68͍!ںT�׀[쾾�+y�c�WY�y���Ŧ�91 ��;I�p��u����~k�z;;��vv_^YqI�*D��v渖�8@�	x�A�<�+�ŋ��� �def2� ��|��o\�B_��s��B~9�6�9�U0"���&����R�JKK�����Lq+�M�-��P�rz���i}o'�:�V��޽{�j~��^�[LRPXX���TU0˪5,��3y1r'�f�=j��/6[�����egn�G�</��F(��wM���4<G�3nh����/ETQB��֭[!s��JX�hhhhET�S�/rr�k�WA�;ja�K�r�q�N�ڕN)`���;��N��$��X@����a���S��{LR�\`�[��'��I�|��r�������^P`���A9�`�N�E�*������=��M%� �@Y�ѥ�C#���Oz=�j� �JKJ��	N3M<<��^`��ÿZf��Õ�%p}��$/o�e�b������~��pFL�V��9��V�"2�x�������<��-���7���QG�slD.�}�c���{�G�`�{c.v)��#Z����	� 3A*��yi�I�ni��'��҇Em�2�e��6�5_-N�dUF� �����N�
[jPɉ�2��$��Px�����oh����Λ��Ȍyyd|P��nP�FG���,ژ$�(�����Q{�V����t��V���!��a1+�z7��t~K���m���0rn�u��8��Ij�ށI}D�A�o����D3�i�y.+?���<��PAk�ï���a��bP�?��}*���nT��n���FP�hm��H��ijgoof�ǂ �,/7@��s���5�Y�11�����5��S�+�=)�Aɲ�,�؛6��BևT��CԖ�~8t�|*��*���w��<o	뀂�6����#���ZZF:o��D)ceuݠ��+�V |]Y�r;$$��퀚���DChe�B�y>�/D�y�����R�4�`�l===�es���S�@�e)"����C�j�&xWy��9�045`k�0(s<YS4�8 D5�ė�.Ng'��{	�.%%��*<��:����+��&ZU!\2d���h�����AZ��WI�1�;�v�f�o��Z�V˯6 �hyO(�zw��:@��a��/��@�q��v+2�[ �CjWv|���iӦO3��Q���1�?8J������:��*Z^t��^D8q��!dɛ7o��w�xf�ޚ���ؘ��j��5Ǫ�!��J����Sn��,_̢�ի�����ѦI 6��e8�}oo�N�Ү-a��t���_��ca�8���	�晱�a������4�}���!A����<��U�Ǳ]]]���y��w��Cy�RqE`����l���36Tg7f����E��l
���&���:  ��ɒ?��2�&�8��!����&۶�d���ا�GS�1��9�L����e��x�H@�u]h����G�N�8�D%��#����.9�v�e>mG|B�Y7<_{Bt��ߒ0�*u����Qq��á��pA�𖰣d��H�C@Q`,Pt���N��h�S�=YN��-$x�V�;��EUf�ΔWuIGb� S�j�F��4��ܒ��]�� ��(U � R�hU͟C[���S��!L��b� ��q��������j4 �N6���7��xt��pE�ޓ���a���C2���J�����n7�<�U���9Z_1�c�����	�PD˜<�-Wn`��g�wP"�8k���O>�jW�h��8��K$�ԏ�߁��sMT��o"���	�$�M���f<�|�\nL�ɱ�b$jNЁ�ˡ�t�9a�ǞT�m�H��i$k~�H�g.��"�4���17n���I6����o>)>�l��͕}��|����x� �ٸ����ɓ1MMM$)��n��|6�t��Q4�D�TA0/�r�'��.Į���_���Cfl�����Ty�A�W~��������0A
P���)�."������"�Vq��h�5����#�\!�����u|Yҏ���j�Wz�]Q�>�8O� �ךʫz�+rk��7���P�t��B^r/#;;{��`�L���S؅��Q��Թ��jXWU�j��{��r����k7�ő8ן��"���&�9��f��N�ɵ�-�[��o��ͨ�NUUH��!1`&�<
c�W�M�$�w���m	nBJ��|}���D��}��7�&�R�b�>DE{zP�/�h:��!����_�Z��"�0��j��7P����c�ջ�ě&j�~�8U�_�;��~�yPґ��J"*�����h^Ӻ�0��@ظCU�HK�s�旹I�I�����>Lz/��F ���X����2(��:	�����@��߼)N4O�Eo�ݸ5��@~d���Y 	�f���w�׶-���G��c �������vm@1{��y���������ܳ+��؇��Xo}���D礏O>�k���ݷ��sM�2_!��T��i���<By낳M:��ও����0�z��Ɔ��`5j�#��
Q��	��m�^�M:@���(�@����h��g�\���K7�) �/�k7߀L���Y�*"��7�rOw/���Q�����=z�TyB����1�oX��L�UW����A##Z�f��9�����G=|�EO��Ɩ��vS���sՄ�g%pi[4�/���G�7w�e�CK�<�ӯD�Gg8
(��*nZ@X{�ӧk�}��\��-��򭪲��s+�ړS*p��J�34�KE��w: a��F�?�a S;~;o��ic?��_<�u0���Eԯ���P?(͛9#,���x�n�V����or|�EDE�5�ֆ�䖏��F	h_R ��C`XYɧϵk�Y�$M��t@/����Zû~�����{m�[,�!��m�UT|heM_VE{qBu�^'h���@{�ln�)-'�-�K!��5=t��ܯ�7;���^VV��rA%tl�U���>E8�<�H܈J�e��r?:�
[C͓(\�/����pՑh�E�cǎ�ŝ�a I?����T�{{�������'x7�����i��"���s�~ϰ����}R0�c Gl�W��a!������tt�[���&�߯�ߺk�44"��)(�����ܝ2!�T�}#��,D��${ X={VZ�7��x�&k�Sc����L}�=y���,��:=��O����_�"�����G"Ztb��\�m�>�>��v��	������!�{řv�mio�!ع���l��n��!��^^������ؽ�1�TT�'G:ϟ;W�ݲ�)�^���~����2�� {���er�~�����a���;O�f�� 1�n��m}���\A[}�^���jD�b5�0�¹h��{AmiF+=f6�21�~���)�����5BY������2ؒ�1$.�#����,����_�:I�^���YR�I{���B"����̽GE�6�~�0o�=8ߐnot^����]n��"H�*V�;\��b�|��)�H��9�"�'z�x�v|������/'��_ru�[������8���F�̇b���S��T(&�K����?��R�r�A�n�H�Y}�/�(�$a��9���4��������[�|D?{�C���q	=���	�{��Hܒ��β,���| G꣥���_*�B�7��⡣�<*��,"hh��ꚱ�Y��@�pf;�ZW�������U�! �%���0�/^Ƥ?4�!c*fz�w���ߎ@�������}
R(�V�j�`Ծ B�	������T8=>�[A���sZ��h��t�^��s�=�D�QȮS��%�T~��t�����lvh ����N9��1n�u������Ӹh}��-3�g:��FۍU��M�.hK�(����KfA��k6m���{�TR�6�up5�����ƢFr�(�(�]'�h��pj�m����h�����bB[,�c�
�9}l�y�_��C��و~� �RA]Ą���ui���?{F�q�tM����;��Ũ+ܶ rm� ����� ��� l��W6SUy�b�\���DZ�Ԑ6p(��d���~N:��0�Ҁ޲!�@f�|�+R�=���A9nbf�긨�T;�,�l����h�
-��"�� �7����K�eP��RQ�8�O�8���%�P)o/�� ��fYk��L݉�*v�`� �����I*��"T	f.s��q^�c9rǒ���+555�ܜn��n��^�z�*Uy7f7?�Rq�J���!m�%PIn�R��U���J��-���Z�I:�]%���ׇ�Z�^���J-��B�,���vK��:դ��Br�X��Y| G��$��&�V�K���
qM.p�]�T�U�����4;���aґv�C�-0X�摦J�!��\�h�D(�F������:Z�0���9w觽x��&r��~��W[�b�o����2�u﬽��t��4���7H3���ٯ����廰��UUؖPƏ���"eCD�*��v���r����e����2x}�/h��.�Cc�aqޕ�GRԚ�8L���s	�dϐ�� ��V�2��IJE][t+����qe%���f���Gϟ??�R�Ә�赳��8z���(�������㼯��@p�S;p;!�^ǬuF�&��˗r�XD�
ѫ W�����]{͑�?ω!<.�*_���I3��͛��O8�"�D����Wo�fgd�}xK�ѿ��F��R�Є�bF9�Gf�NMѪ{Ƕ �u+)>����`�˃kײ賴O��M��A5��1t�
,����!"J���ns�9��ȱk!D?s&)<2�ulBh���+�G�H>k����[3��X���f&G28k��,�e�.���5�7]�te%�$�ț�^�ƾ� /��l����f��u J��1�@!���Rc3Z��X�/�k������h�n(��]%����}��>М+9>�| ���n�FFF��p�W���k��q-�5�����YSW�ìA�b�@��~�Q-777��b�L���\�Rm����&���Bs6*v������9yF,T�P'Uq����O���yN:8��NKk�g�
��lW�G���՘5��E򷬣,������ds[�������0����1��o��u�H�߽��_���̌H�}��{	^/�ι�np��nh�|�������O�P�cA]袣0b�׈م��
V���4�\�~����X�R�P��<��Im��>�N�"���^C�~hh��3��d��W��:�}�x�kjD]��l�;9w����.��@��?c�回�6�Β���Z=������ΤAȠ��TwBu��Y�.���4���q�Gi{� Ru~���H�I��������伯�ܼ�ҝG5�T>�놠�+?�R�]���艶h�$� �G�j�D���40Te_�3&}�o�N%�_!>�Wg��F{���br����K6���}��ᶗ�԰P��U�B��~(��5����'6±�7����!�AE�^e���t�*�j��K@hؿ����F�cd�4��Pd9	|�
a��x}�ا�*� �1��TBOeU���6oMj�O  }��e�S%A4pd�Q�΁t�ݮ�ڥ�EpC�ѿ��ű�5���?{$~s`5�ǐ��c�v�8��:�R�����jjR�{e�n�47��S|��%%y�����^5j���܎F��p����S*Z���[���;��zC��v����*�Le�c�u��iiκ���S�~����wTF�
>=�����D�}O�O����m^\�v���0�3wwE
�����P�Uh��܇׳ڐ���־Ҕn�V�3x��ܷ��g��c��C��4UN?�s���]G.�?��_6��n��`�B�}O 9��qR��V�dR}/*E'Ɛ�J�J�4�����	��<�_�'�f�G~��G�����O�F�m�F �j�Z�&�m
@(X7A�Ъ�l��J���egO��`&�ܜO��!�z�B�ugU4"��h�TV,i��QL2����Ǥ]�}}}jّ�
-�䢢$�=s�cI��%����J�sݛU����J}>v�)��pA�1�y]���I�rJ3=}���=�J6�t��ܓ����3����'�!�%`lz�����D����a���!@���ґ���&��0A��Bp�ÎSo?�f�))��F�� C��{A"0�u�E���P��/��	�Ѵ��׀�| d�|�[�Q񻼊v\j|�Ύ�s��!	��ϲ�P)�N�c0�5K�`�HDP�����|(��s�9c���WN��y%���J�$�����"�*/AD|M�j�w�7j������ݞ����b�L�l6"���:�	�%#Z�����(�0�U�F���0����~]�믐�cц6�^�4 8��J�Y	�b ٝ��F���e��&��X��4	��sKJ�p[/��,�K�v�p��C{�^��� ѽ�G;&cI��ٞ�`Cc㻸x?ת�mnh��BIՄU�J��r�B݌���L�^:A ���c�|�}�x�f��S�����;p_�S������|�q����+��+z{{�~��Zm��R�~�:���˴�C�8�Iq��T��<6��'�_B&�4ѻ #c�i]��0��ћ�g�R�A�R(�X��yK㊐���ʢ@T%Q#������TG��,�M`������F��K������L}� ��bFf�Dϩ��|�ѿ�鞆FN�9�R�H�$�`K>��?Fی@l��#�9d�ƿ�7���=G���Ǐ���������{�5�c@�<��gɂ�htt�$O����<fiIbef7�+��=�i��'ܸ��F x' ��F��ы��_�� �βqla��Z������g5\	�8S���*�;�C��ܹs@{�Z����/ßf�O<�!������@�zL�ihBj,������z���&{�%���|�L�R¾צ�	~� �T�
Ϩ����od�K8w �vA�TY�4k��E��!p[��s'.dc�4�,(�Κ���|VA��/��+;-[�hA+���z�hÓ]����m"��fblg]�D�^� w}�����0��;}a�z��ϳ��qwڑҳ�����!jN�3�PE_��=��k�gG#�b�-���z�kc��WY
_u�����AAA�"5���P��\j-Z\��ڀrЙ��C��/ӆ��m�W~���v�+���b�jh�O�hK�r�Y����V��R	b%_�j>��F��ޔ�~��y�.�<���������Fp�n�h3"w�=���4#bu�U������N4O*D;5�{��x��̓J�����?��}��l��l�*l�
�zH�	�� ��k�r����d|��1�^�tx��%K|�A^u�B�������m>�	���&��
��]�̻�Zlm*������}�ݝ������Ƣ�SR��@kL���%X�M'���/�	2��J_��`��-Մl�ŶV�<n��,�FЂ�S����6��J�W�0"���'~�BnBKW�ᯁ�~����⤻����N��~�X(��w�A�H��@��ƶ@�啖������$��b�T�`ccc(z��5rD9-/�2%99���E�sá<4�]a�h\��m��S�hΒ�lE퀐�����yF�' ��Y����t�N3�9�'""�r�Kx⡄�goo)�~��>f���<KIYq���1��d��c���������+W�`/�'%�]�@\8�y�1���AMӱd� n�قj\��L�� ���YH�����T��7M�362��CVvG]̶��k7��"�(i��~a-=������x��OO�[��0�? ��V�\��MY��C�b����$D��p��8��卙]@���{���t}�{�x��g��B,
�8/��rBv��G��'ћ�t���� �(ĳ���_y#^Keu��qSX�9��;�c��*�h1
e�r�X���#���)�!�j����df�l56~����c?���?��#j���H'���ߤ��P}J�B���Y�VP.v�v��,�1��|t&lEG�ӡY��w!z�Y_�V��;T��i�o���BuXS����ڏ���Q�`�H�=%5U2,�Qo��Bk;򗍛	D'�@�N%����vq�Xj��nVR[{�Gj�a2���(�������ǡ�N����7fـK�߿ע��-5E4ƙ�*�Vnz�Po���x=�3����,�첲2x�-.����eo�R@����2
�+Κ�)����bxr�K:N���ڕ�� �����������mS�{�ҕ�d����Ay,������O�Fu�eg�-��Eo!��\QQ!��e�W�Pg�q�����;-a//��o+Z���xN&7�>�}X ���S̲ɰ����h<ݾ!#�̘�VԈ_��t�{�N����GR�JC}g:0�#.���UmoAס���9�����C�H+)n]����w���&�;v�y���v�G gd��3�ց/��l�������z�n�T�P%��`�'M-�C��@�r�[u���3�Bښ������L�����%�#��cA ����M��\��qIQ)K�JHʾ��5%elQY&k�d�:�V�5{�qJH��K���S�X��${�����t����>ק��4��������y�!��R�m�	�~h��:|���A�rj�S�T^7.����˫M�-���a� �O�2K�"v����7F�t~�D�	^�P}?x�16��!��My�_��,���{(%�!Uy]s����#�������4z��`z��	t|�l�c[1����w�L�u����Q~Փ�"�.`��a�aA�0m�;EZ�^Ye�^2�hy�S`�2��}n;���X��1�����������{@��q@��ՌZ��B�i�J�W�3���yf[�>e�]S{���ֲ�[�ڨHr��In�{><lq��L�e���}<q����,���\A�E�_\!���Ӆ���;�t|��@t�I���_!Q-XC����o�ޤj���^�-
e2����Ѯ�3��$�c˳��͛(�d�e�=��p���iYY���R�;v@͍�d��O�ty��k=�ȶ��>�a��	�cJJ�kݕ�	��O|Eb�������g$��)�W�
c���!�� �Z�x1����א��'9*�;��wB��*� ���	;�s���I5�y���u�6/�m����M�峗��Ⱥ�5�r'555|���e�R��?�Y�^^F&&&Z��NbO��2�V*A����03��e���|��v�LB{�.��j7ev�  �_P��e�9,a���vv��i�t�g�t�������2�&e[�-�pq�������ϟxh��~K�ī"_�8v�������%ܴv�q�}���RS?��|���V����!(�pA]��9�/J@�aԡ����B�'���H
p7������H���P~�KK�TX�lon���?�	��ڋ�����gDq ���m���w~�(�����`]�jWր�nq��^�C�,���T�]�ꏱpǉp�	�.���sߜf���p�Z�]�b7�A$Wj2,rt ��Asm�گ?�]Y�ɇ�����[�tx[����}�P��x����"Cu�
[l��E6�ɌUo��=��,)5�:���
�F$ ���:����Õ#��?s������Q�3ä~�'Z�o�%a�w����^�D��;�-��H6��1)�Z��nD�l�;wP����=<�>�~�W9=�r�I&�����iA��P[p��g]����	��i��3�R�p��E��>ii���Smh��A
~��8����J��SN����}�/¡���5:3sV���и_u��­9��bI��3���+�8���Z9�E��fX)�����;����եw��?����Q���v�}�k�.p��U��)�t{������m>��?�6.�E�'Ϋ1D�y$���2��w�#MM_|��M���!��#OY}�$q��b+���A�"�M膖���e���t~�6�&4��M4�g��U����jx�θ(u�Ν���P\K�ƹb�����h�"��<9[� 8˵�C**�yyyOJ�GG�=�_��5�`��t��<VY��u>��ǌ�v��\oooQ}�<�����<fnm=�1<VYX8˥���xSw�[�n�B �E��=/UT[ۡ���L��������ϒqA�\��@Kծ�]�7�m��Pɡ���Іk���mmzzz��m'�R���-藣��̰�%��߶� �l,��^��G�
���"�%���F�����KݓySQ�˥A^_��yS-ls�@��EQ$
�%@�F��.h����[h�G-E]5�X�uS�m�Q�`�S�1cQ7�;ޯZ�n:r�*;�yG3D���	h�}]ޔc,�1 P��K�ɐ��b����3�<��[m������Q�����.Ղ�/���M78�����ߢ�1�$EG��z�@�@>�f��Ǆ����Nn���X��MCGggۗ/O�9i�Yo��C:����11�(䡽H�E
tq�LL璲˷Q���U_�}�xۇ��m�.0B�����T'�w�0�6�Җ�s����G�kfv�&%m�Li�>w��h�S�����CX�7�!�q���,�O�?rn��I���mm�2qC"��r�/��a�,��ꁯ��5��&31� go�Um<�l�dõ�k�]�r�g�$�d��l���`w�EBh���@��t�u�Gߡ��+Eee��R�u&|��O�5�C�O'���f|AoBd���	ཚ�W+e �j
��ΫNsUT�����3;,g�J�\
������EQ�*hb�cUr�Y%9���}���t�AX����E����׌q����`�|6���+[ގ�_��!�
3]=�I���,��Ȁb��q��Vp;�����J�]f��b�>�AV��|��e�FK�����*�3�C��ki��b��}��qk<詚T����Z������}���`��T$CX�y��b!'/��}��۷3Pڣ+�^���bQט�mѻJ�y6��I�>'''2\#ഭ@�\E���m1�Z�~�j�)��a�8��鐽��'�?ߝ�:=�f X*Z�$Q� 
��:�"e�o��Wm0�R��U�Ob<���~/�@�pCu]� ��#١�+�
f�#�E��D8ޔ����
���@�Q�?**//��xs���V��e+���5i�y�5۷o�����׾}{]jz:�n�ά����Ύ�#fU��:YZO�zj!�`���Ǐgj�ӏ����[TW'��%
Ԫ��ؤ�.��MP�y0j&���R�d2�^ۦ�ΐ�T��	z��E��p�ތlId������p�(�v<&&F�):갾CP�E�r��K״�[�cd�.,�U���� �v�[�N1qS@�<�ua�����+{���g�ѧ���/f%J�2��m�g�%��"D��LLM��d��Ǻ�@���t��>�ˊ��X?��c�@9�"��S,s���|�M�@l�舆K�Ū���� 3��_B�����.���>hd�w���������:w��������i�9t(j+*̅��&{�|�<M.�o��z�e��A�p����;�6��b���V[���dFu�\�̭�,&�jp����S�H���Y 'p�f��o�P�˗�8ݱ��D�P���NL��kuva�P��D"�����e/���D�����N?`�B�i��$�F����8ArQuu����g��9�R�6mz�5�KT'^�3(H����b��;�Ah����>��Jc����t�(����9�qu�ӧO�ǡ�m�0�A���i�%���R� %�/���*��uw'��$g'(܀ܣ�
�M��m����6�$����x�!D��������q����	\ �͛[��a��vӉoA�f]�&�ŀ��,�R(�ѹi�U�u$i�c��OB���Ԉο�~'�rN3����Rca����e0����h��!����Q�ﺈ_C'�=i���>K���w���Έ�K�����L|�����}%K��뎎��?%~�Ӊ�韯=����ǿ��Kv��+���:�op0y&��b:��Z홐�8�K���e^7?��ć�"6?��ުz`��������@��Ʈ"ss�8�F�Ul-s[�*�!���Xyzn�c��09v�)r�U//[�h��C������pH�fT���"�+x�4��C/0�p\�+�nFo^�����^����=�7箩<N|��nu'��)l�V�%�����;QUTZ���	�E:�v�ny� Hft��))�\ܔ7�}�;�W�'�_>�%�<d��ȼn	u��ϟ>_��	~�����Ç�WJ�6g�W����lP�s
��K�켪!�j{�S���Θ�0�h�ߥ�!�S�P_���H�m���3���6u��`M�1�4��[����������a�o+�����s�L����P˲ �ݨsK�v}I���pŜ>�6��c��������n�d�~���w�-CfZ��;���a���������5.-I:Ar�$:jnnT�_6E��4���Ҳ��9�o�:P^��,{���򃈽���7~T�9?/F9;|��^���^�ADz�{�IX�F��6 Xݨ [N<QQQAV�)�����8%� �0 �*U�^>�θ~�r/�n��O�-d����p����btQ����mހ�@�B*	��m�����)c\�w�b"�����TH=XiM{e�t"�x̂n�������� +#��[u�����5�Vch������b�Z��zmDJ =1��e����Ր	�!�"z��@,�<Y�ZFb1��ja�?R�:_Qv��AV�>4�
�'�@�dj�G�b6w�/�2�<��D�UW��׎�i���ީ*<L4>��(�����o5��uT����p����Բ�[_K�$D򖭄�U���<i(��-Snn������l�~�1��J���f��a���o�����)h����P����ȿA�����ā���\�&���ג0C�.(,ܾ�R7�gb=B"\�(�5��=���+��k�6	�-���S?������&sD��_��<)=��*�`�C ���KBo�_�AA�?��*����N����#�u!��S������[��T�L�'񤣏K;�(�߲����C��M�	��-�}�� 8���}�W.H%E��V�v1�"�:��;����W���B��B���O�CU�u�R��
�k�'ؙ({�lw��h�1�Bᶧ�/�Tx_��z���*������7\<���XA�1z�?������dDe��~2B(�{�A�"�
}h��B������E;����~;|���l��!U%%��މS5uլD�w^�fU��j�_/�Y���)�D>�YUC�X s[ ���CQIvySV��
C�z)n:��"tp`����4/Ar�玿w:Rғ���������c�X��Zk��@U��gq�@���{hf��,��E2PΠET�ٲe�ȷo->=-�i��lM��H�F��N�����^���
�.��.�%�~��g~�R�ˍ'����ޓ3nt�t�*��;F���Is�;���W_��A���0ILcZ��AAveh� ju�O��D؋/Z޾��)�}�p�B`��)#i��l7j�LN�\��:A��Z�s�<ٜ�b*<:�d+�V���S�}%���04��H���v}X�s���pV��hL=�� p�3|��� �`$Lʩ������Th�l@D���b:��th�P�'��JN�6c)tS1��^!�ϫ��/ΗO�.����"3s���g�!uV�C���h)���USCƸ�UUФ��c ��K0rX	���o��:S�{(�h�j�g��DFF���u�۽�*�����g��|��Cvn��WV�����g�rc�!���1#\����r|�89�d��˭�y���E���h�
�=b~�WNEf�ޟQ5$� sB�Fn�Ǧg=-mEzh
��E�4C�� �C��I2����*���2���$�yۼ*o��PYع���\��> �����W��D�� ���qC�12��Vr1�����Z�t �;�P �R�Ml���@2�EN!4��~�m6+�-v)�t�G9��3�Hwv1�ؒ�L��2���;��n��!C)�$����7aa��K\�I�S x*'�.mIv���g�c�w��8Q7�0��,�D7�B����������~�"�g�6b���	�@�� Y�td�3e��d��d����5�r]H����f��O���7�\<���y�Һ��I��E`�R��w��E��̦)R`]�l
���в�XK�19���t�.ߩ��$1�D1�p[�SF��I�.�f&X�Oh�'��BF������>�[��C��$�p��|��	fɿ�{zzV���(�]�6D����I�3�r�{I壣�6�ɦ2B��N�-�_�t��+���y�5�Jǥ6��\��H%,9�ə������~ͯ���;]�6�X�^���Ѣq>��e˫��]�M�茞؃ѫ�P
�P�� �j���$� ��Yyk��w�\m�zt8�I�4#�8��.���\�N����I`²�2��>�%k7D]*� ��G+�PK���^��!�pN&S�+��.�'{�_�jlU��L}:3��`�4��ji���1�ӿL*n���)��.f��6(S�G҂����qbFVb|V־��������}Y���U���:�7���-�u1�l�����Z� ӪU�K���}��;1���G0�g�4�,g8���J�g�w�/��o��x�~9&h<MU����G2�YC�.�0�c/ЩW�����!W�f�d4�����cV6ciiia��D��G�8�q�_���䝜��K�F���[� �<�~���+Ҹ͇�dEDK�D��&wM������$E�e0C%H*���_6��^~qg���a��ɛ7o����g�R7���O���Np��1=��f2+�����װ4�3��� NPH 4~�����r ��^��sLC#������k�Hl��w��w�^�j�Ї���a���T�Z�����Q&�n���(��Jd!�cG���.v�A6�ə��j��.��;@K������z��v��ϴ�3��$�j��נ��z�(آ�"Ѳ���u��v|�u7qX�����z�C9݀��T�C��l������ûS�8w�2kim�G9�Q�?,8���Ը۷׹��4���~����:n{�Ϣ�G�jQ<f�����P�`a/�LBC�\�Z೛D�їM�۝�C#b�)̯,����L2Vn�B��WL�� 	���c�����\�_��}j ���l/��[]Y�8�5<s��&�2)�L&b�
����{���~�j���Ӥ߿��y1�o��,��P����71 ��'"[�r(�?/'�r(-uؽ{wnccc(���ʌ����{���{ƼWǰ� S�F��7�ZzY�P��������2t��」fC��"���N��n�l���]����ig��Fՙt��m]{�c�L���n������#k�N�鋯Y+��j�V"��8����:�$�F���w�Kz�%��;̆Xwvv*u,o�a�\)}����un��,�AyÒ	r�:E�gT��zG�*�w��w�d���T�v�؍������&y�P|~���Z�n�?kP`U0�%��1MRlm���^>#��u�����:T���Q��[f�+�r)�I����@�/�H�j�i=>�2���Y�F=�e���g/f��0;���L�8gcK٤9O.0K�O�?���W��4��������5�O��+*z=�� ;�:��������![,C�	J�Z��a��U�h cn���b4��@5@ä9U�۶?�k���Z���`�+��5O�jTx�L��^�;�w1�}�=N���t595��;�oJ��ttj�-�k��9�[�i�����w!.L��s�Z�v�~��Xj�ܠ���%��s)>�T,T����R%��I���4�Β�zex�K����R
E*B�)_����XC:�A�׈d�7#�e�۷�y|Y�,���ˌ�Dh.�n7SSK��܄�MM��=�٦�e��p�1�BDӥs����~.�	���$=̓���gD�ӵ�*[����^e�xN���]n��B�6��en�ii	�3F�����������JTgo`xY��;"Ld����-,-S;w�Z�FJ��������~~�.���T{u������1εp2�3)��2����3�l�'��e}��뎨��WCy@�-��w#w��.+^F^>��!PVY����eo��0wH�G���u����s��r�"�
�.//�È��~1�$z�μ�>��s��1�<���i���M^EnAU��D<�?��eww��
�h��z_�8�##'��2>��%F-������fl�UÜc�l�̗�f��2�KAsV��I��ܓ<w��6sKK���44}1Z;������322�[�[�tA�]��^�f�iF.W�5�:V��w3:;L.*.ދm _�x���= �\�*7����O4��N�� ɝ���Y��q���][�� #�<������K���σ�ysG�s[V��r�?�q6�ĸq��H�<���_��N��-7��)jY��>׫��= `b����� z@}y�� ����m�f{��Rpx�T�E{��P�MR�U%�#�F0�L��/)�sHEC���\Y�V�I�Nk�t�L��d�i�Y�kgM����~:��B
��)��8��ɛ���PH%��;��SߜS�ֿ����	��	5?�S,p�$7�8nѻ���	I�h�F�Of����1)t��kҰ��N�9���k�T���<��K2�n��h*ıu�ge�޻��v*~[s!��Ȼ��E���:�:ׄ��G�!��H_�rAlll�AL����j͓�e��(Š�A�c����EO�m\����4��)�uܸ�g�;��>Hs�*#f;_��N'ϜKv���3��/�x|M��p�ܗ�M��
�k�����ѤĔ��������Wp΁h6�R��ك\_	Dd��q���W���j�R�i��0��"
�l5��|q8��{n�����}��͓G�����䍻'��ů���u��y���������CZ���(}QJ�R�V�O���9�����ﳐ���Ѵ	C��.��Oh�v%(p��"Hq�
����zV��$VV�5�CA�v�,$�7���:�����Ѵ�ꁣ������,?+�'��P�r�����WY���@���/�Fv��27�L���j��v�c;3R�Iz@��|==��c��а㪟���ˏ����8���¿E2����܄�q{�X����a��΢߿~��X0�`O�)H�K��~�ɝX,#�h?�V����L�mN@���p؁=����v�v�T�4c�����!2�,���X��+c�[�Pn��G���|?�Z/��t����8:9��tP޴��h��
z�6g����'(E/&@��b(sh ��FmY��mMn=��#ﮔ���pɿ�k-s�2�0�{5 �2D�=٣K����	��M���Y�Td�̖\�a�hr��=ep�ر�G���~LM����{�����l�`� �y����	"r�N|?�Y�8��c��/#�$W*�_�m�;=��S���$�ʹ?��ў@��k����P|r$�$���KHEI��<.!�o�W�ou4(��\"��U�/
��WR V;88ܦ�)cL-;F�F�n��^4/���(f���X6���������4\�rhF�$��@��n:�o|�`��+�Ru�ik�㍟f��G6�"�fbz�k*�����i�B�Ą��hHk���^Eee�J��(hh�����x���Ȼ��f�[u��B�����>he��{�wl�ؚ�'�Yņ���^0 �Bj�)��m���Q�2//#4r�a�ӕ즫N#���!~���M��˿�KP2�<�B��Jݣ�t�K�� �����f[S~߮d��� v�X��K�y�#�=��}��D��{���"��/��M*)�J��v	���Ivv'(�",�7lk^�_�N��J&�>�Z��$��_Q�bA�I�W�l�W��x������U����u��u�&W����.Ɖ_�Q9v��0�ˡ�O4CZ���X�߶��\�ꁗ�.�"�)��yɅ��us(�o�fԝϻ��k�cUS�
z��1�f�$5�==/uo����	����v�}|<+�ͪ9R�O���[Y[�k��f됈�N ��VV�?<�p
����27��'7&��.�����δM�z=9l&�(��x�c��'����Z�Nn����0i���ׯ�$�#s1��o2�{�MG��0�P��S�G�����|l+ҋ���E�8 2�ӟ̑��5�u�32K� �]
�mHI�źs}r�W�0T�ռ�I�C׼&�qh�8;[�cz:���t�l�^n\�67[����oh�d��"�!N��@���_]8���&�����T$*��a�BX�8V���,��B��Y�X;������Z�6�5n�m����E/���pwW�	��$�m��{mw04y����K$6^����M[����w��fB��P�,��q�4'Ԥi�U�Do�>p��v���P��~273��Sxߡ��ο��+P�9����!uUh��!`6D���?��~Y�q�h�F*Q��Ka���ɐ\e�ph??�h���}�8�y�8@�da��G
����0�}Q�3�S'T%����D��ʢ~�|b!PG3�#�?/i�B�@���h�fy�%j����
$˴?��h[�ǩ��FT#ğ>KnG%����-��X��S$Y�^���+Ի��P�L4�=@6G3��� FP��2{X�U}hǿ�����)�3�j˟�"݅�h7���ssGA���<�*�OQ҉W���^�STX��9E����T'����<��ğ�0i���6j����������9�'S��QZ>/��� �9p��)�	D��!�ݜS#ny�W�u��0�fI �5{	�����<�wt`]M$ذ��lܡ��A�� H��a�����c1��P����_��d"��ı֟?Kn�J -����^ԍ�"j����	�ի�U�#�q��1C�>T��o�����SiQ��G}s��x� $q�RX,cw �1�mL��������3k�����#{�AԎ%G+Ŭ6�ѭ�Q���+��1l�"����m��(gS���Ő��l�ǎ��N=2�}����^~�'uN�@�رT@�	�h1��Qh�tmva�Y-��=whz{����L�(6j��i��q舽Um��2{���Lc���t�.F}j����؏��
P#s!�_�B�|�F��_�:R��r:,���[�Ti������i�dkk�	q�tү��J�N`j�8'j��SF��^�S튜�S��c�@���p	3D�"�h�R�m� �5'±����v	��2��W�`ћ���H�Ygg����h��$/y����z��R�[��;�@4\�������4^�yq�;�Q�Բt�K�2q��ܛ��]�v��]�t!?:�p���-��y)��U��M`}��i�%K�����ݵ��1%�����u����h�>al��cć&cz}�f�p�I	��:�W/���������e;���c�D��l��JC���Qޭ=)p�n��9�>-�yT;�/�2�R6)nķ,�ŧx���Z�_3��RF|ts��������z�i��`issū�Z�(t(%b���^UYƒ�2����wg�
Qw*T�v���[ڳ�<y�dr�WuC
�m�-	��� �Ӛ�R7�
�2feeV�v̰:�I�T'76����B3T�g���\��c�������-y$Î�yh�XX[�Ƌ��2KB�i*t���p0O�*�.��%͝u�~q_bo�u������q�CC�d������u[�.s���1A��o+�`����xm��`IEE�l�L�c�$�J����W����O�x&�b�����?M�N�׉�*�J���3��G��e������k��Y�LF�D��̦D�>��]���%=�Iae��[1�*�<������@�ȥ�!Z������� x ؾ>��E{�Ņ��8I��:>=Nqx���`�)�q=xvM�e�e2y��>O��L������?�*�j+�E���Uy]Cпx�d�e:zkH4�yì ��nqY�C��R$
���^�݁I9��6mB��N��u�B9���&]�3뼔q,^��ʹ.�"�yX)f�jo�s����q�&y������?+����xF�*�@�(��
�f�̬��ē�Ca]��?����CS+�S�AN�N��~)�#f8�|�'lq7�\Df���e����Ɩ"ֲWJEz�Z��Q�`3l����#����ₜ܇&�U(��B���<��D$���_ȩ�����fY_�r�B����P7
� D�
%�}����h���Qh��OFȯo������LLLF>��|Q���P�y�qvѯ�-�:g�2���;TQ���U�3K��)���XV�.[o�T���U���w�6Z���5ۿ�m���b��`ͯ��G�Ï�f����#�Fխ�W�	�}x]�$(k�dDgg:�����`3k�V�WA�=��_5��;8��/��A���`��кF���s��X�y9��x�M�ё��-A�5��ZA��
-J�ȵx=�oK4V��R����^+�}�e�i��hz�����މ�j;nO]�xq8z*"\�_a!��AN{��Ƹ��Q|o{�����`q;����%7	x�܋�tz��!1IX�6�f�}���$S�8@N���=��i�S��V.��Pq_���:H�۷���O@:%--msjr߂Eq�8~TQ����4d����Gp��C����x��S��j�<jҩ�C9Z� ������/�����o~�q�� m�O�4E���Єk9T��/�[�~�s��?f�T��r��W�{��&]l�@{&q0o����2�u���Aǫ~��q���w�'���VWW#�@��Z4k�۱��A�-�F>��0�
 (����_���q�Lڗ���Ek������+���E�F��GWC�d��"�xrD����4�����ѻ�E`i�̊c1�U5�J�xJqF�E�1������g>�(�'�^]���_�.�yR��bc��MOT�YL�,�(�S���/��]�P?���m�h����k���
�����v�9�2ơ���������
�z+Kѻ����8���>�i���yr����2?KB��v_q��մ� ��I��i��YvM00ff�A�ir�����3��z4���5���lİQ� (���*�Fjݼ�6f����4>�T|�=ʥ=�ekd�J3x�U��hc��mf��']dS��!��4,���ۮ
���z�N�y\���yU祜O���h?�W����i�h�eX\��8���zl�+�:b�ò��fQ���� �WVJ.��0�\�jolE���Xl�js�R�ǂ��+>�Si��1�bu�k!'��߾M�=�d9���G���MvF�ˢ>�R^N�
��Ц��jҾ����qwr��}�(	�Cǖ?^�eH\Qln�T���x�&���ݽmv���0�S�+=���v����v?�Х�I�#c շGX�/5X��5��iXXE�0���@�v 2vii�N@1?K����(4���x��K�o
?�����KQ��zҤR����2�|�ӆO���Щn�O����J�����.���ؚ.j��P���}B�>_��X���g��?�qddd|�(�Vu��:��8�dT=����m\\��,,>��[z��[��v�MSd9��\,y_�ް �S���1h��g�Zs�8�˱M����6pT�=�;H���V {��O�"�ɿD ��yu�6����?���]$�����B�r�:͗;e��z��b$PS�5����w{hu%��6��i��X�k���<�X���U�(�q_D�/U���8I@�Ᏽ�r�޵�����紹�{�M���J�E�����:��Xj{}ɚ�c��GS��χO�=�=闞�����k"��?��@H��T��Y���q�mW�T����y�U
-���Qnl��l�ws#�
p���.v�tJ�c��!���IF���۟$�y6����M�L\�|��Ea�9�k� l3���f?
i�������Q���y*�R���7����R暵Y���� �i4u�կ3s�fɿ�|̴�ᩰ��:��ֱ��k�lͤ�ß�� #�k�V�=+1�0��q]��~V�r*j߉��7���ky3�ZZT�$%%�HNHs�=Z�'� K���'��)��z{��с�D�w�=��R�!z�����Fv��+�W��ʐ�:�e�ն�vJJ���x\�k�u"��'p���+\�+����(�aԳ����+�T��F���b���0z�Ə8��"V:
���n��C���l'�5,����	})
J��̖G[�6#vs��3�%8b������v��!$�2M7�˼����X�2t�ʾ�&�ڸ&-�!�k>���wa��
�(b�
V���6
K�.n!�<p�Nz�3	���i~�{�́}J<4�6d�ӑ�V{�P�_�<5�J`-�=��5�ɜ�_�<ئ�.��|���m�x�W��DB���99�X�&Y/O�!���.	z��~w(��`F�pZ�QØ����J^"��p�'���q��Gr��P񞆒�����_ߨ�|xN�?�X7��B������G�3nd��傪�v]E��pӧ;����/�i1�`f@y������k�D� �%��~;�̟Xy�#�L�)���!oQڷZ� û�S�{��ԉ������YVH��{x���s���%�� Ԗ�<�t{�M�3l٫y�`�1�ϩ�������޿��H\1��H��Oַv��K߹s���I\I]=��;�!��y��,��G���P�jfww�F^bD�
;��[��h��c�፟�7�8����II��ҥx}!� �a���������= E{s�Gع����!�%�U�p$(��ӵV��C\Az�6n(g����7�z��	�FNTa4�UO�m��:�ې}��7_�^�*m��y�9vߞ@H�=p�L�:�<vѣ�sɑ3�=���A���/��Ï9��QF���y ���g�G5,?����7笄D���f-�
���J��M͟���]	)6�߁f9E��(z�0�����Ĳ�����ӎ�~�)�������w�$�l�Z�n���*��G.��g�& M0�H���N��Ț�i�\~[�|Xē]+�  ����.z[���E�*� �����2ν�� ����֒�a��L�Z��B�2�
��@񱘽��A� O�X�y0����.t����v7��f����س<-�.�bB�wԶxʱM���G�\pY&�{�o�"k����ܼ.�:��v����}�p��u�3f�'^9�ץ�C��{�ee�����Ž�mjkvb�k#z�)���!V�M�a�z�@��0���g�gO	� >}�$�̄X�v�m�Y=8t�M���)�H���ʒ�բ�R�i@W�L������N�����3��i a�p�خ�$���v�yS�a���g�V�$Nr�+/w��=��N�5��m�B���+�B��O=N�yK�y��(L�K�M�/sB������a�++u���er�p۪<	oX��L��z�M��p��vXT�]�^�6G�~}0h����s�]�����>�ǌ�_��.�Vi4f�Z_��1�
��9n�-wb��錃���))2���ucܗ�
1��@�4y	2=H��G6�gp
���i	��7^glkw
���3��NV�n���ʤ�u�B�K��N����9Z#���g�KT�"��Pf)���A7Aޯ�=ASR��^`Y�M?L	0g��;|l�?�]x�`P��<�s�O$ ��gĀp�5]�e��`��ڼ~m�А"����E��#+}d�����ǘQ�z%��P\��r�U#L俕��bz���0D��/|�Ty
�}����������g&���f��S�+9��n���;اq�F85�Z�j�q:!Z����1�9��Z�;����{����6�Np$%ef�./wz��|�g})(����Щ e��=�`�G�v�����	3>N�f��^ġD����T�3T4�_�Rk� ��I_�զwt��"�?q(�:㌪P
A'� ��E�lS��z=��2i�k����a��P�
�y��!�^��PYw�Nj�bt���􎩩��@[b���e^�2�A��@�u3ͻ<�%�i��nLa'@0��������a���g(�`<	�.�o��:���d�׳�u$���4s��u�ͨ1s��T�:���ݻ{�F��;������>o�|��(�I�i�:EhYo�k������jo��p���z�4�a9��G���׎�z~L�5䍢*�6�?��X��a��m�uu���O�e�3h�0ve�M"+����:��>MSg��5x:�]��v!��{�n�x�����W�Tp�xlJ)�q�m��S��L)����wC�F +}��+�f���
�wh���s�k��9��`�6F��;(��.n#��=����C�	������`�j_�l0��:ES��h,$<�~�N#f��g�j��p0�+��O�T��c�e�nA��!F`�)r��l��Oc������{��ۋ^��^�8����KfFu����r���wy�v�e^�e�]R���(4|�m�E�ѷ��A5d��!9_z"X������X�y����ʓ��d/-�B3= &]�N�雯�}�n@�'���`QFTߩ[�Np�{�4 L��WL*��{���yrr�XJZ����Z���D��c���R��`b��W�'�?{.I�����7�~�ʉd��^��=5ϋ�Bn����x,?��m*@������M*5sqP�ʤ��a{0����S^y=�j�%�/�E���1V�տ�س���W�^]O-$�c��ߓЊ�x��q��<�ÿ��6�EH���+��r����I�sR\�����0�[c����N��ŋ|��{�j,�d,Ve!Wܭ�	B䈓T��c��w��o!
Zs�gE<O��T˔� ֓Sޙ�e%�i*�لvn��ǓiF������ r���䞗�at-�z	'9A��!��Ke9.ԡ׬<�A��wU���A��s7��V(C�+�Ǡ�%��OF�r�*��83Ѽ�H��XV�� N?WC��"U9	Ĳ�t�G�K��q�"-H3���s���E5�6���OB�SRR�	��ΐ��G{>  ��-6�=�Ù��Bm�Xz���z0fk�� �q����r�j�6��r�v< �2����Z�w�>@�b�WВ�侣a�R� �gFߦ�:��:%�5tz����|_��.,���K�F-�������i1�#33�"�d��-˿@���+�+�k��_g�}�_iW�sG��f+�v̿b6-�.��r[�S٦��ZAM��}L�(��6e����YJr��z�S��� A�����X)��먠��J]�cG���S}7�_��ŀ���T�!��������=ZV���ݱSSO�5h�Th��U�3�ÿZ��BM�f�N���������G�m��ۏӶ���;�n���7��&��+�P�Y<�f�B��N�����p:��<Bz���w�\Ȼ݃�9׃9I]a�T�)�-�0p���|+����+Z���D�QNV���}�?��#���te�u�A��g�,]�����p�`T��v�keت�~H��|�
65̮;@�:��g����zy����0B���V��Yˑϻ��O�k�<iwt��+�/3��חL�hٛd&st�E}����~<Pb���%%ig���t}��!���X�9��Rh��"ע���
��ChWy�����e;]�����nՔTzhw�֊�2^1�3�zj|ff��Ӂ�Y�����r)_�<�t,V�P��[�,Xj�qܘ-��TZ	�y��Ӝ��@�� �"���%P���>l����T��{�����z���+����Ӧ�gh���/Z<w�F������r]�Ph�=��b�U�zX����wƊ�N;ǣ��^�{%|4���s	�!�l
z*�� ,22��!�$�(�̖�_��%r�N�Aʿҍ8b����;�����5J������7ꧩ�NB�Hr�=8����Q��j<�ֿD[�,�C�,�u�6����./��D�:�UV��� �V��=���h�"V�����3�-�r�mA���h%HI4�	�����߅�3з���I�}tg��A+4������]�{�MCw��;�&��@�����S3[�O���W+eT=�����#���Z`��� ��V��a/4ڨyT����}h��2:�h��3:�m*a��ևV�}�q�F>��?�UQ�KN�f2�]�a�����{��֦h�ń=��J_��/��ս����$M�����N�J����\dP��<��������9���w'����h����<�W����3B�uXZx�c���2�m�Rr�~C����<,����ٗ��� �w��/��^*Y��e��8`�=-��n$���r��q�y��(g�� ��q��L:�����ۨY۳�A����Ʒ��y�k^��s��P��/~�>O�Ĵ�T����T�S�(y���En���>��xjy��nQ��h�5�� ,�KjF�$��'�!yڰ��P�*O=�79<�u���X%���@n6�{٦���UD�4Zx�C�����ا����_�<�u2b�ݯzh��+���3�Ә��Dz�1�s����ron���;����n�o�=��W[Q�l;??_{�Xǈ��7�	n�jZ��h��ڶ�T�P����6�=1þG_�u�"XY�l�`0z�!�������OwA�z�?&�:��2'_���b*�*�*�ga�zz��������"x\��H�I������cU���K]�͡8]*�!�|;�B5v�gp�2�3�nn����Qu%�Tnm{k�����J�)�H�
!�2g�<�SH(2e:%9��y�2%ӑ��<��M���w����u}_�*{�k=����������y��� �M��~���3L#��8�Gh�Ժ�^>u0��hyrU�W6ve����Lh�ڧ΋�2���$h���d���ƶ��F��y�V �.��XO�{L����y��������v������o�3D^y��{&�ڐݝ|D�7.�����?�{z�w��w��H���{��|�����4v�=��;���6+�S
��/�(�v���Q>��N*�2do_�7�O��REj;�g{��R�{:���nn������u �~܋��B��L�N���)ʹ�߿ӊ@=�[3_Ih@��czz�����6�j� �ȿ����x<EYl'n�3�n��8����|��J�ӣ��G��U���s7so%��X����@
�_-Y��c',������D�:��ܡ"MO�N���UCv�������8�%]��$zN�fS�M��0���:�8���q-����n���~_;ww��65���~_&JԶ��z[6>� ����?��M�*�K�&����D�Md��L�Ulkn?�k�Q*{ӌ���i�{��x���{'i��)y]�HZ��b���ʱ$���G�~;��l��:@�;;��5ǘ�d"�� �2۾(�̰A� 4_n��*�>i�{�e�<���.V���KS�c��I�����"V�=<�G��LĮ���ԇk��DT�����@f#���k��Ag��x��aMu�^�ou�E���qt`�O����=�=��:/E�����~sx��P��yapԗͨF��`c֧x��?F'x�>ǿln����g)�\([�~z�馨����-�LL'^G�x�+��{+ȯ�]��.�z4��,�]|gI��H؏#�AD)�u��-<�凩a��w���8P#�C�p,���|�p%�!޸@;!7V����.�T�ǡҝ<��_�%��z�/��j�'n�:�K�c�G	��gc�_�0�u�4�]xŹy�C����[s����Sz�Oz��%N#���#��G�W=�|�*���^t-���=f�s��(��`f����/�{�����(w��Vδ`hM�'xC\�ja>{n�nW'� B���=�7��J/Ǿ�a��&߲?E�c�������V)���5��KY&�Uӎ�#�gy����EK���^��xL����sT�Ǔ=��E��ru���DP��)m#��f�#F�	=�����i����%y(g*x�o\<`j��j���F���F!�+��>����d>
�f��
}#�Ī�������E^����\.�a�980H=C�P�=zf�%po=�D������G�mvڄ�f��ٲ��!Ҥ�ݝ	<�U���~��2�0�%3����L��d�wk�^n�炷��
��9����z(O������ �����{�K7D�V��[o��s���/+�U�����P�u[	o�X��m�#�-5d�%�yz�,5Vi#PE&�M.���f�**|"��E�"��3t�����o<L���pX]i	�Gɀ��F�×��|��|���</�P�FJS�R���G��?�Pz���kl����޻�{����kY�@ݏK�� ��Qij�CK�3��%R!��w����,=�ZYɃ�$ɓ�۷@CDL�~�[�pt�b[����)m3v��o|�Z9Ϻ�7��������踙[Z�r���@E���2��{�k��Eh��z�V�]C���PWgJ�6��[Vw6��E>��8sP�P���h�	�x��[*�O��v�cc��z'S��@���Vs��~:�@�5u��'Yrx�拨��l�_��?�ڽ�nq��("L؉qV�m� ��{�(x�2��c��N�����6��ǻ:G~���?O[`\�����]��7������T͔��)���8�m�Q��(
ն�,G�s�Y�R�A/��p�FaR|��p'����;��٨��{`ew'M���&c�u������e %�ݍ88Л���r�x��)��������G�]��4|��,:d�zRh@iK�ݍ]��c.q$#1�Nr��as�d�fJ�v��Xo�h3�)l��Eb����q��B�_S�]]#��S�����#_���E�����	0Ϳ'n�4Yꋡ�����ϰ�FOj�o����W��8�4۪k�is(���7YH�v�e�?a1ů�R��+o1��<����Y �{---�}}Ǣ��8�TN 8^ZG�ot�I�	�����g��0���M26���24��I�K�h���g�t��P��)�Q���Dﬞr\���or8��5��F�l�j�9^��y1�k�=&)Rn�z�hʶ�ҏZ7��(*�y���"Q�}H�'�2�/�I�DI��y��6�=�Ex��9�C���QZd�qzl�MFq3�t��-c�E���)9�hn��6��*�-7���j���'��I��
(/Q}*V�����,�8�����""D
^�����%}�ZdV�%��5/�J�T���ÄV��*�	�ҔgMMM^,�bt[�� ���L��CHՠ������V�@n��2��Bw�<����
N(��X<|O�9.����Sa*���|2뒀����thۑpYa���8����:��tN�XZ^�$�Dע�!67]�h�*d2�X��5�-�{��QG$͖
��7�3�uD#�`��p�9Ξy��'��@{[[++k�쬈В� c�r���g���l��X�����i��ƥB
n�1����Li+-��8�(Q����-N�CC0(gi�f=�1A`���Ĕ���F-�{z�}D v ��a�m�� �LK����fs%��=��h���*�W�������Ъ�y�t�r��`�1ћN�}�fe=AD�m��Ԗ	$�+E꿃+���
QI䂹|�� !�>�|:7m�]̺{M��$�aU՛�v���z��[�9RI��ݝ�s��uw������/e�����������b�p<���J�)��" �|��φ7P���<U�ځm�������,7�!q�/#m�Y+�-$����rk}�n�ĩ�����?�t;|8����. d�	ֶHl�H�v"3#�~Jӧ��fvu���O�����Ig#��4�ݪ�N�j�g�Тk�[�L3	�� �8����Nqq�}���(c\n�����잨!��:���h�}�d�O�#��ш�d@^]�q2�U�y�0=9���kL뉟_� ���qn��ǺWw|��N�C�>hV���Y%�+�ɼ	�h���>+����p>�:�R����jѝ�A�|�^���bIv�,=�ZL[���~�z��W9/��p���	��B����T������?{��� � ;n�n{0�y�F�&L>�QDvm��҄8A?�*[�̗6��������Uc�5؏"6-:�-���V�I*�G']�AV�8�G�;=;�Oo��zf��y�P�N�q��6���������v��4���$C�v��3*ɏ��af�#_�V����k���2Q����_V�)�QNJE��GB����;F�L��4�ۙ������nݕ���FC�g/����r"v�k��l���39�����S�ȯ�����q]��g ����e[ngh߂b�NbH�d|�A���S�U�'"g*��#�.�#�����lO�:��y�=3/�#���.�41ISK�Kp�"�O�1L��m%��F����(>Z�9���E�NNN�<��|��ѵ� <��!W��̨{	���;�V����	�t���*�s]�8����r"�z�n�}+6����	��`$[����S���W�����%?�_sA�Ho�+{�R\��tZ�˖1n$�<�����π)�U�#�����@:��ȁ�j�cu��Һɷ,s�����Cј�])��I�lT�Z�9F�s��N3�P~~��9~��⁵�L�L~�=YU�)� ����?w����Δpխ��	1�"vB�!���������O��r1�:v�1�#�Gښ)�H�NO�lc|@�d�ܯE��g���K�"���A\-� ��Skto��g<��^�}����|��/sVZ��g�߿�����fV�V����ąȩ���������_c�N3d�	v\���L��Pі4��ΠS�t+�Q���#�3~|�Գq���uAn�$�f�:w�vJSHl,{fnn��S����S���eh��h�^�M2;�^�OhLr��hw������>e1gSs�T���=4����Z�F���7�г�9�inZ���i+yhL·�+2����I���
��lX��م�s���w��)��R��H|����p�ʂ��S@���z��gH��^�W2۾�6p��Gi������CA��κu�N*�ܭQe,g/	2���4ƥ�f��o�Ϲb'a��@Z.�8��N�/
�4P�W��9�illl_Iɓ�&�����$�NJ��'�����/
./,�Q�;As'5f����uX��t��I�/7l|��y�*��qB�C���(���񔮔<�&U9��U��t�y�vᲛ��eYjn%)&�ra�	��v�fP���!o��W�O�m�f~.��~���8��I����m�����)���z���C�:W#25���$Xe0c��D�����Pw��D��������gZ�Q�l9=�}&����w,��V��5o%�b���n���e�<Y5�?ZQ5dR%=�a��zN=��+ �GM��=����Q���sn�ٷ3\�=6yH�Sx��s��h���d�.�F�ß��a[�fI�x�Szݍꨠܻ���1sHռi��ƴ�S��]-(�A;	�4p��g�Ϳ6���my~�L�Ӄ� ��|ȗ��ӖO�%L�ݽꡯ ��C��>(���y&j�5���Zzh���FK�^���zMII���^�e��e:���7�98>)&�SS<�����XQ�&1P��w`�	C�*��L��$DHd���k�tήT<�"c	IS�6tus�!O�]���EM��ots{"Qot*8�u�n���tW���8����9l4���Gw}�LI6��Ie�\�7ꇘ��)'5�z ��|=D�����>]jp\2��+��4���>��t�ʟ~���*t�{��
������}#�3�d
�Q��lPV��V)�:�-�S�M����-��U��_��o7f��|9�f�9�,MJ%�R�l�/���rb�&�xv�T��Pe]�CHf���z�)����]n爾�P��C����I�(��(�"���"dK��Yr�W\�gf�7M8�&�Bȼד�DJX�z.�·���z�<����e;ry*J��L�f�i;�4�so��fi�9���a���hW��ӕ��ŉ��+G@+8���1��f	��%��WGM�J���s�?�	ypF"�kw��1y*ͽ���ٶi�k|'�,�A�a�����m�-51'�KD�ڍ �ʏ�Γ�؁����L^����k���0���.�7pi�q������d(��>{ۮ�#�~l�t; ��xh�P(m��q��+��Y@P��#0'�p�>�%�5�f-h�:���+쉨�>�4�X"E,8�\c���\f?NA�z#N��o�Ҡuwpv�<\��I�C����ױ�{�Bs�h6��o��e��C��ɷ�G���ft[V��:��E
�oQZh�w��F�S�[
��#b8c&�{����Z��S��Aw+�.|@�P�]j�[dAV\� �y?��GZ�S����&�ZQ�x>��3D��U�=��=�� �����j2����>p9Z%�\��p0�<K#��S!eeb�;&�AU�s@�rk�ro������_*i���o�i/�[�C�S��n�kY��݆�	R���=�-�H�>b��"[�n��Z�T��.ۚn���&4ƣڪs����C����z\��Et__l+�z�Ll�w1P�PE ����޻o�@82 �EK�@� 57��M��]<p�P���n��c�ج#��<��� Z��2|�Z3�\P[ppp9i�K����hh]��@/r'Nw�wJ�x��A�����h%쐩�)v��pK�� �*��gf_��f:]�{!ߚAj��gW0�X a}2�L����=-�)����������d�k�_i>���};���u"���ENNfx���d�A,���Q���ޜ�u^�@OdL���g�F>R�<���s�ι:)�1�F1ei:76\�^>pa��Gwqt��훯%�e��&�n8	��Q/��awF>���w�k���r�

��C��a�ٖ��膔��v�$�t�aF|��Ds����tg��˘�Nn�Ԑ�6HCg�_���In?�s	��L\�H�D �r�ne����k�+..P:�R�ۤz�x��_((��h'��Kl�eb�]TP�L�
����+X�S�Z�W/8J��:uA��V6�\$d��Sk��x�5Q#�/(�-]\���:J������L�!^-�0ǟ�
�v�|F�,I�i��v���⪍8��@�3Q5��NwŠv�M�f�1��9�V�R���� �~i�ɹ��YU)G�u�n�U�uvg�_E��tS��"O�w̥a�f"�PK:Zu�L�` ���^��Ք&�Itg���o�'��%B��Nkc7(n� {tq��V�o��8u �\��w���.����S���O��u0C���&Sg[�5���o}��p�Q��!�]�6�B��kS�;���S����\W��%����񬉉�tA��7�d�z��O�Z-�Ln).rG�I��BTO��^�SI��9n�/z1�k�(�M75���;�>��q�G�`ZV�9���^m;t���N���Jc|��y�%q��M��ih����*�b�7:I�{��|40@��Q#�g�
v�?��$`-���5�ӠI�{��&	��n����V�>��5P؃�0��0aƨ�3@CYHbb"�'}I�=�<��WC��pF�����.9C���tcA�}.N-�|^����>�		��lb��rv�	c%��3L痥oH�jvU�6�}��i�+�kǨ��l��O,�Go���>JCx<���8���g��ɼl:�z@7{��g��o����9Ҡ�+�Ɉ߫s>��aI��(yϴg{��}\���I'���N�ԋ�c���N�>��B��h����	�5̈ܬal���zt�����n�����j^�:![�$�.����l�����������ch��)m�b�I���Xkʰ5�1�����E��A��^Bb�o��|��B��y��&];2��|<P��9�}�N
��0?��;2�������8Փ�� ��� ��%������U��O����e����i�=?b4��\���^�S�=���<v�3��kf�\����JbTvS�v���T<��� c*^"������r�$��-`�u��K�+13��k߱@�� ́T@�$c�\�(mMS=�-WOmϳ�גϣ�$&1f�A��?��ްtT�e~�x+:.>�4�a��,7|}�g�JCڄ�!�%#��Hbr��
��U+�r}�G@9Gǂ�4� xm�h���:���̌�������}��Q����Vm�Y]3yX����3�X���|�}{^��\MILm	[ݾ��5%zn�i�o��}��ܵ�RX�ufGA(���H����5��!�`�x��=��[,���d�ch�"�� ��wY�� �)�/��yM��2��Y���_s+�H:��vؔ]SS�|�8ݙ��e�|i��Eʗ�̛Xl;W�[�����Պ����h+'%'�i�ńi���rVL��%���6�`>{�l���y)���������e�/"I�c�,��G���������l9�A�=a����n�r���{���3�1I�$I=�P�����-H~�ƣ���i03�s����F�-��=)M�z���p���4���(��S����˩����j�4}��"q�_Ces�����PD�����gdC4�۝צ��D�%�+�G����/�3��E�
T5��<c�?�����P_&�Y�	����M�F���
z�������Ӹv���I��� ����2t�c���>k�\Nh��1)�CW���r������ 	=7� z8�������~p�����WB�Ys�۬��,2.�>��$TA�xB���������[�$#GGG}�"m�D�h�LEŚ��*��1_�E���[Rc���3�c���_�6}n0}0d'AT�(�WSCѮ�0�p�q�48����nb�NN����ʆVV����z�S4S��?�{�R� �斏 �L�å����k��==� �x��z������q�a��r/Z�Oƪ�����lm��m��tt<��2q'��O��8	m�`b�F���{���K{Q�A2�{(S=���
�m/a�&43o����o9��N��]��#��w'2�P!�[.�c���mȗN�"���߿���!\�k������r{�����+��T�q�݁�I� �n2��>3���|�����g�lo��>V,}x�T�\���|�\��5#c��&&�q�	n�x��JFC
����D�������|�]�z��(,,���dΧ�!�u��\^�o�Xm�1�a��s�@FiǍSa�"�Pm�R�[̖KA��uuu]�ip�=�f	�MD� z����r�M�<|������q;.쯨�XklkLʄQ��/,���ǭB��벂>�����V�<����/ ���Yۖ��Ⱦ�K>}+¦��"̴sq�*��}K3�%S'���͛i߶μ���"/uX'tL���C�O��_0�J�xF M�ͤ�a�ޡ���̶���ãy��B{;::�ʴt��&㫉�U��]�]��K��3�w��}��]�L�R�ڧ"�����4y���C�@����1d;���x<��P��h�b}��9��A����5Q�5Qg��$���099��ߥ��]7�a�{�X�8(v��޻�;�F���]�J��ܨ�r,��*�Z������������{��Ԅ�#ɿ7��Xa�y�%� �q\9䟖	D�����s-�͛.�i�v�E��o3��R�~:�}�==T�ɓ'�W�+��s��x�Q�V�lʜF5���O�3��<��
���N��&�BuM��[h����?ۋ^���+6uw�V������p���@%��?�'5ȫr%d�i+��/##�a�d�ˆ�N0B)�����5��!�P�{Z}�ZC�]N���H��y&+��~�	��?~D�rr[�{�N�rj �����Zc�������d���� L#���(��m~�/久pg��[��NCR�����Y��B���)�o�t�v�1��)����6��+%�2�!�Z&���(\SU}��*�h���";��V���������t?� ���� p�Z���.^?���"��fzv�ET'LL�˹��:q����,����w��}��޷��<K�ΤjNhy�gh�]&���iD���FT:���e//��(�#lx�e����������񱱵?��Cq�;V�=~���H�p8�	�Tf�C����'l��rܗ�@&j�Ͼ(7�nĉ?��P*q�`��#dP$095u9�I��;}�G3{��Q{��y�m`H�KdH�`��>�W�xC�����s(�ٗ'l�
(G2c���\��Y7uw�c����RG��a�&��b��fP��+y�	���="22����M����X�{�M��8���B��{FG�|�}�P�zWw�0��r�7j{��J8�Vl{����HK��qqA��ښ�A�q3��0ZXXd|�r ),x��#�_
����b�R(r�l(I ���<���(����Z(��ʍ�Ok��ځr�]=�v�������υ�m��~��"`@b���{���Ǌ�����O��dFEEEFEU�/������C����X����I���K����L�����3*w�g��~dh�%K���J�:9���� �n�'���ė�z�BS1�	-F�wn}<هF�o�J�w������y�D3��{����?�9
_���vO��[Yc����3i/�kjT�QB�'8"�ۛ�"_�:�o�݁��$���&T�YH��/X�"���}o'3����a��
��`9CN�Tӝ��+�����_�����z����;d Rhi) $`��%�����˂���[�w�+����V��sUm����4��aی��W9kr}c��^M9�:����D�L�w�dn%j��AB,��BR ?�q���|4C~�6Z�0��̀�"^�f����Bo���`*jhn~
t!z��������U( ����O:םo�&5�q��v[�P�,��k� '�żc�4������Cn��ܫ���#��Jѷ��� i�g³��ӕ�Ӄ~*n�ɑId�S�\�ʽ����$W��_��zyOETC�ж'@)Fp�r�I�99���n{ �h�Gf��Utm���C�ܢ,��>��q�o�w���/��綳)픟68��n��Lv>�,8x09�@%0��TM~�*�"4�����k�w����-=*O��d���b��+�L�7�����ݖ&G���}�I��H�Z����9��Z�=�hoh�����=�~r\�?�C�1}�
�w����X���44,���;�1[�	�C�|n	�H0䒪�j��5�D����Ba*�[�[&H����.�;w�P��j����菪QDN�t���' ��އ�
`�U>~����O=:9Ay �����ւ����ԌJa�m����F�X�*������udW	��
V�{���kjk/��չ������΂ܱn'vY��MEDaڂ#�a #߾}QEd�,m�Un=�|�pm��f���;�#�^olieU������e`���>��"𳧻Q4P3eQeazo:��Lŧ��Q�Uh!�����_�J���ijialIu���f5�X��6[	�}�1�m�6.(��&0Y<��8��v(�
�-����H�G�vvgP���N��tg��l*��clsI冨��v�.�ѯ���.K4�622�
����e�c��!//��g�anO���j7277�Wx�� ��_���ѣӌ���&�P&�Q�8����X��l:4t`R�4ac���b��̤��;�������V�l���������W�T�Ԇev㺡)�G=vVV8m�L�9��F�xy���ϰM�u��RXϵ��so�dl4��M�W�>�s$#�0^���I<5�q�z���_��Y)���̶��m7g73ڐ����9[�ƙc�Gp<���_�����xH�p\�'�
q��7~�JH)7!��^E�f�C�����Z_c�5���A&Ofֿ�!v2�yV�DCp�)�?O�~ѵ2�0�2�K���'G�^���2A?U	��b�A��qT	�	����ge�C�-�<���h�,�	  ..��Ǆֻ�q3�a�C7jdi�++ܣ�q�<�_Q����3��,�������L�e��l�P��i�z����8_D�#���Zc�YWk�8�:\P�F�!p�	��#%n�)ɇp����uu�0C`�FΌ2o;Վ�N����|k�>��jZ �B-0(㔣�H"�\dɱ}
�rc��(����	D@��n�N�\7���ŉh��@��r_���;oУU��Vwǔ��${D7�7�	H+�RKOuUJ����CΓ����R@�|q:�<Ɨ���ٖb�9�7�g���QZ~@)��L��;��X�u�`�v@睝�'��A����������mmo��E���p�b���:�+cI���,���f�\p�T̌~v~���J	b�Y?���6�� ��T��Q�6�k��[#�h��7���wy�
F ���@��t`�s<�]!�P�@1���]�.p�6��;��͗܎S�D�r�ރ����h�H'~������������u������A��+��E�y������v�*���@{�e�����LS�裞`��Lu55�D�*7F\����"=���]C����ԗ�����]|9�%�?���7*��ª�½D"A��ރN�Q�H݆z
3�O��,�Dp݁c�\���+��U�(���P�g��1ۤePƯ��	�{�bi6�N�(,H>��J��f+?�H}��!�9�p�=Ϗ���j$�l�2�_�f����:P7��\�܆4������B�����d�1סe �:LhaoMo$/�P����>�������$��u?�!�zp���p;�H�%�6
�T\Iu"��皙jizm��Tn�j�[qb���j{�V�.b#������~�-w�s�j��
������w�9�#�E�]@˵ƍ�;���s�T�R?t�c��Z=(��]L��{����@HPS�?�xa�n%� X�ݖ�;s65��&&&f熪�ra+7R�3lM�v�E��;�(ή���%5�>sƑ�+**��[|��
��pjh�1۪���� ZgQ�ƾ����rp��3��x6K����f����x�	K�� S�1`���-�Tէ}ɯ؏SP@�m���l8������^иQ�-�"���R�$QD��2XnUO/��USZ�Oȸ.������#����E�(��[�`ڨ�P>��>-F�Ipxd$��*x?n�����Y�ZS�[��$/�y�w<k�+ww��a�?xQ ��(�_�L�w�^��}@���{	�mjjB"��<����Y�ڪ��>i��`�-���s7��:4#v��Q�#.O����ʈ��1O��#�R�b���$�痢����k��o�b�$P�m� �o����`)5�̈������_rs��Yw/�?��"�T�sM���x'����������Ւj"x�_��4Μυ�X�O���v�e�4���:8�C�A`�l��F�쁔��trk�����Dzz���0�z�E��/�.��rC�"	z�=������ &T�y;��_��P���:�����e\�����,N��n���SpEK�8Y���$�����.���3s+����K��"48_]3؋?~|Fj�Q	f_\��$�B�D��;ղ���<�YK?��aF��Q��&�=�j�bI�t/��;(À�'���տJ,�V���
y�A�s����������N���0�\=JS|(wը��s9r�F�'Tt���6��gDΟgDN(\(�:Ѝ4���ލ}/�箢"���ڀ��V
g#P���9E}�>�=�s�����>�b_i����ϯ`8���/��ˌ���`�)�w!�j���إS
��1�UL�#Kf��nt���e@CL�0;�F�)W�E9)TC����}���Cc-8��ڋ���tJŪ���(��;7��ӛ����'�<T�Y�Բ��&���*�xΈ��
�1������A�fR]�{�� ,lܳ�wu249f��.�[p�vе��$�ɬ�k��n��)p]ktZ���m�!����h]��YI��ט}s��,�2�8�7�Y��MKR�R�]�n�r��V�Hs�@��=�H3E�h.��L��><�f���[\�|�-A �y��,���q/�sf$��~�Mξ>M���P2�'М�����������y�b��C�[��^]��w�K��s�$�_��2Ϗ�ͬomp�.�z���2��3�겓��k���=�����A,m��~-���W�Fxp�J-h+�1�����I)hA�赁�X���<�F��x��ɓ�it�i��s�x��l�?H��(�U���̝��+��������8��tv
�l)���X��}�_tr�7O�qq�ؖ����A��4��8���q��o����׾�#�s��k6�L�=�f���	��x���h,;]hG�Z��eu�Pey S�fJ���$�%?�Z�b���1���2����~��Pn��t��Uk�@J���X:Nž��/��Jk-�]��~̬�՞k��a���o���=^`�-M�`DC�h���*�G�ҽ�'Fߢ�w���K%�Ŷ��Gvj!�O�ǣ��S
��m�0�`�@�	�}�Ik�ϗ��)EK���n�e��^܌.�!�
0� ��d�$��/��<����#��#�JI���������D�.0vh}�9#��I\o�AD�ꦒ'�YS�@�7��gQ_� ��.@�~D=n?�������J�~��x�,G5
���A~	��H�U
L�ag��!m��"q�,�+fh��	�9��A6�ve��ϟ?+�?�^[D�Q�����2�8�t�_+M�P?������m�2�j�E�G@e�:�#�e��h��y�l�,"r���S�0�M}��3b�")�D�Y��S�Fk�h�պ��IB���U@?�o?�.�5�m�k�+�P?���k��lђV����m�/ZΠ�w&m9��f�o2Ƕ�ű��/�E���D�w�Z�R�ȪS��z>�|t�.��6ې���C�|�)��5Qg�Rff&�@##ٻ���U�{s&4� 0�(�1��r(N΋#::}�5��O���C��ѡMkd�����Hٔa����CD�oHP�K��H����ƊVJ:����]�	BNS|V+�����k&12n瑯��AB5��@Ã~����z�n����z�qf�rvى�L���"���y[��rdll t"��7� ��6c��323C��G/3��8��{�~�֕�Z���J	~����9��O3�S���Ͽ��m��X�m7ڃ��X�G�̱R�G��v\�\>C�@#P^^>JZŠ$��k��\�Xa�)}�T�58ྈf�d+떖���\��f�V��$@l�KW���G��hI>|#�֟�
 �8��=VD�Bۍ�a�g͔�^�1��(�m����/�oa�m�m��l����yQr�	�t�6�~?�n$:��&^��O�}�	l�����:Ց���%XJ3^A���30,�iR��	fv�Zܽס!�((`��P�)��>�����$�^k�h5�b�C�����!`����mv�8z��TP2�C��8R ^W>��e3��*T��4�鯖��魅����S����)K��(�^��P�L���Fd���Y���[���Ds��L/���.M���a� �񒠽++t#�N1�%��>Y�d�V��@�T��eV��p7��nʦ���O�_���k[��� &�~9ʀ\?�*�W�(I'���H�~�/�����A��.��xl�bѫ}�6�^��9��h����u%�a8ۺ'h}��kVؘ�s�E%����A3e3J� Yt�ћ�E܀�z�1U�V��8e_"�`@��� �K	��_%Q5rU�^��	}+Rq��y�@(�-:'��bdY���R�fZC$�F�̃�WzS����� ;$��J���*��Fo���ۊ�fMD���P��OaO4tqȺ3C�QtF>���m?����� )��2�
T��n�%X�R�@�3�8�Z�hY���.�ʹ9;�B�Pq�7�3��9�w������U�^wcT_0bs�l7���PY�o�ƚ��:,��I�(��D����K����Ef���O��{"V���gB���l�؋$z��A�О$t�E���f���*o�( *��&��I�7&r(���8�����J��`���������4|9��?%׉�+�~*P��9;X�6�ѭ�pi#ss�Q셠k����#2�};t�Q(z4!��J7#�@_�/���Ӵ��p�?
�.�����u6JNk������ �y�	���ի�ɽ/aw��G�"�{<Y���1a���WL�G{��+vgZe�������*�o�3|���k/�3�h��&A�2D�Ñ�l[�����$��WE����Awp˸B�[�<˅v��­,����<Q@�.$�p�6�IB����"���0|��,8w&4	<��<£��0���K��X��c���B�Q]�sz������q@#��L;�� N�T��1T�pc���h&���0�$��lZYg�ޭ���0@���`T������+�X���D�}`n�����/(7ZD}<���nT��X��vF�$��&?~,O}�7����7�T�d���ޗN]k����k˓����ԫI@J�� ���@�1���	� t�
y ��cok�o�4Q���G3�7ʺ��ܤ��V���w%�i9�'��QF����KCW���Ǉa�d��D۔!�w�7��wJ�/<�^щ�ζd����E�m,�6
��7F=7髦��b���@܅**1�R�Ƹ��e�����c��J��@UC�R&~�rS���n��]Y&l_�C��]Bve4�� �#o �`>�l��š��03c3�&��MD/�244�ZQޗ�����
�I�Q����-~�,Z�C>4������]��BVt���uh�04h�r�N���N�S����!��?@C��+�;�����+r��J��\؎�J&���B:��h0�`Nǣ�����9�M�DΝ;�%�W�,�2�%��X�wb1����<қ���`T)`�]]u0D^���A������$�[���f,��(O��J*ڃޔ�;��ʊ��� �Q�p�n��ܠ2��`x0�)�)r�,r.�&�nA� ��ab+m�.vL��;�h�sZZ�NN�-iwΚ��B/É����5��U�q�jx1J _FGb��т	�e�㑿�7�~�߈c��E,��;���}�N	PTTT��Z�_t�Ooj��^2֙<sF�5�e�L�L2��ENs;��pw�����ԣ(��--��{�7�q`"E�W�Y�r��!�;	�(*��r���HW����זa���0VD9γ��@���ѱN�����]�P�c���[��W�-`^�?A��g']���<r>�𨪺�^,���`��uP��A(�+7?�È����0��ê��q!�F���p-iU��̒g���A�y��`WQK��)�� -�|��~]\�c>;"Yp�l8ۙOh��;(�<"��Zo�8L^4��������De� #���Zl�6~@�� �hϣ������vN�J ���3�����4�a�xs��D��(�`��g�~ʭ�*	%,V���y�&��<T`�ѮP||0R�T� ԇb�x�=HII�mH�������*�u ��Elha�th��sPST�P���E���8:u�E��Y��aT�F]H=��^o� ��ާ��;?���N�y_JkAC[ h�?��gKvr�u��0��c
<��؟?fAܘz}(h�8Zio�2��)`.А��;g� T���H͡eD+ШD�齂N\�0@�"� �E�:��U)�.H3R���D�����56�\P��g6&�����V?�ۢ�w�@⌌�C��P ÇH�-�8�Ld�R�6F4S�?��ox����p�����f�kc����������C�2)�@=r�+�y��䵏�S��r׊o�4�����wc�Eߟ�*�v� ����՛�eM}}O����'[�Y/�0�������&s����E/Ʊ��VF˷`��������y&/�E�UX�NLL��S�ȿuj=>�w���Y~�Yu�K��f�q���\[_���EA����݅JU�NE^qN-i�Ҋ����Ȳ:���H�6�'j��RYzb7w��cL������宋�.l����ω��dZ��c�U����ʻ������wf�����!��n�[I^9M�w?}��t��^_��5����z�Ћ8H����f�ݻGxV�YV������..���iسaǰӭ��챇_o8�x����b�O��ʵި$>}l������)�%�߰I9���fǤ�{�=��r�(�X��M..N���^����)�RA�;v�8?8�/���߷�ޢs�oA)�}���)�,����.\u�+��pt\�Q�����l��_�Uq�'"�ٓ���)�"�(�7�'�/�Vl�֍�����
febd����ڊ\��7�p���#�z�W�n�J�[j�0Xɭ��&�fc]��j�pqƆ����!�{KKK���d�|�2s�P_���΋s���055}(�޷�G.lp���ؽX�4�䩃��500��f��N�>��ꡎ��5��_�]f���~mT�8|p~�Zr��C�������o�/�b{0�I��>G�k�0-g7�#:+���U�D�J��!����GF}�ju��ċ��u���v�����kF����n�Q�_2�\��&����␫�i��:9������MHI��Z�r��0p�j_��Ծ+v76;���{���Ij��g��W�����$O���5��
ꩬ�W� ��u�
P/�]�
�c���"�������o~k��K��n�-�$����o���D����t����Ф���&�,��a:xa��ę��%O~�'�`ns�~��~X�aF���	*p�Jb��nLn���SV������&:Y-�A��A�z��m������ݝ;wVF���i_���Ż�/wn��'�:��7��')o{��R�Ͱ�:�ô��e�]ң
7�|9)�z��8ne}.A��؅�&�<;�X_��vd�j��~Z�X��ߺ7�w{��������~���#R� �T��E��/�`����X����T0��C��{�����϶Q�7�Z����	���|b�TZ��O�f+�!��Ɨ�eb!�?�/N��xZ蹯����4��컰ї�������

M�#�,�D��Vo\7�\6���Zy)��m#�M{����ڇ.{���;�Su9��u�7�N����������[3���&>�LX�v[Cߏ�z^��S\l�SU0b����`�l�'�͐/H�	yԣ�,..�N��b���gJ�9Q�qA�֒�t�J����=A���o�]�{P���;�(��xM�ל�����QgM��>���5�?񝸀���##1L���v�Pr$v�+l���a�R,��4��-�������S����7�U�$]�9{��go�c�j*u��n�؋�<1����K�����P*�9��H�ߏG��j1�/@ڜN(��8�q@�@~R�W����������r��^S���P������?1�
��&��2X�8۽��vo�ݔ�l�F����ʇ.�T��s�e������k���7�����-
�F\s��֟�Cپo��3���^KHM�R�(�e�P	�$eˮ�죒�V������I�b,%$k	S��l��3���������yK����<��~�y�w����ҫ,�_s����^_�4�G���#徱�O��'ﲾ�K�!Mx�"��߷�D7En����o�ѐ�*�1P���@�*Qݎ��"��Y�D�X-M/�t� =�ssPY����\��������XO���_r�N���T��,�iv�<�P{.j��CO�����0�����6�y����6������a%��TMi����n�+��!Bp�ul`e[���Gn#�ߐ�_	tq|/�0/��6�yA@���?t����k�v,�� �쭭�t�{c��A'h���+�����b7�w*x74<�M��7&��dR���)����%Z�d���Ϙ	��P�+��}RM	�G~TVv�먮�Aݎ��K"�J��UG
ۏ`s#�6Ľ���;�=��_Hޟ�`f��|K�������2��bB���hpc2�19�HA@@@��� �K���L�K���c�	q�}��P��W*��9`�Rw�Pn
��������^X��꿳�[��UZ�#�3��"=�~ȧv��A﫡�oߊ-S<������~Wv�-�<��G*I?��n:$'���lUSs�O"��۳����1|Ev�O���mZ:�,�1��C�&z8�Ŗ��'���7����'b����(Q��7,g��+x̳t�]��`pc�U������{S���ް6M,'�/,dx3�P�sb�N���"вRP��`�]7���m�[�e��LhL�(��WN�	���1����+߼=�]��JVH�V�Y7'�����_}kpC�7����6rk�	��1ֻ����'�	�+\C�>\����L�	j��DM�s�����
��a�꟔�4���8Fs1A"�ߒRx�R!�_�~X.7<��iV����(Xyw�@�t:�R����r�M�����Muԏ�J~Ք΃����ׄİvC���t9v����Qq?�_��
ݒ�9TGp�tl����oB�X?��'+=�����(���^�>�����aF����+\���ka��b�;�o����֖�"�ʎ�X��{]T��^�'_Pn�7���/xa��r�]��%Z�iiK�;n�	p��mݺ��0~➭ U�'0L}{��y�,�İ��������U�|�cN������xZ�Y%A\��e��&�:f�#�`�|�ɯ`3=�Buը���?�GJ�U��xA�u+���J��@M���V�������T���U��!]�����Smh�`x%,��K�}���|�R�V�v�nk���yp��U"���n��肕�g�AJe�l�����*��}o��g�����Ư��g���Tr��'�A�.�'�5Q�9�[v��ښ���O�=�����=�v�y2�7�]R�sq�L7�1�J<�,���$WK���������Pm��9��1ڦ�^�9F&�����:�j�!�J����m�;����Q���+vVK�<�Z�p?Vf�������t��.��i�5dd��s�-��Haͺzz�BBBv�H[S��K嬕�nf,��_���{)BdGGG��ؘ_A���D�_y\~���s��cK���T��X&DvZnL	t#vq�|��dhXX.Wx$���3��������t?��������1ע�����l����8Ḱ������)��8�s����j�5���
�Z�3	A�ao�#�K��QCb �(�k�94E���X�7��-]�Q�+��բ�JQ�~�ѓ�H�׭t�6bC�s.���c���Գ���-�(-���J6����d��1#X2&8z����.ثn�Å�d=�>h��&��zN_M|�����P^̡���")n�����2�x�pՄ�!�ګۆ󩪩҉.��3����7��F���(�y)�͘1t\�c�I���S�|�qq<q		�Z�BZ��ҽ׭�/��G���i�v���	7К�0e%%_Q׃/B���>�l���=p��jFUD�݌�Us�|��+�����_:�I���X�M�^�\:����	���ַ�]���#��`(�֐�r���{�/�e���T�k�ช>ܸ�K	|.���۾�^�KD\��m���=A��)���������7ov�֏�L���?�aR�!��\���h��R���Z[���D��ڠ�4r�=��m ��אj��xUY�O��![76����B�p�෗�gf�ǓVl������8��e�ܞ����X���:\ʙc��
�+w�|�{x,5��9�J�
���֞@yH1ݣ��x��A'.�Wܷ7�j��� ����d�����5e@��^��~��@\����[&�]�x��4�V˯�9�!2Yvq�����v�Ct;��`�&�m���H-�������W+���988���/�k�ψJ{�.T��6\����K$��i�m����#mgl�5#+���<��iR���c`��)\Q��M�~�2r����s�߿;��߉�8ߩ�e[b�Sʂ�6P{���Gy��a�Nrck�ث�i���	�۶@�K����u�D�T�d�c�� /�d����?��4W9�3�F��
o��~�{\���N$��p<%Ҡs����9UGUl���[`�oC�	�^�x����x�ӃƻKI�KI��k�t@�F��
����>���?�F��u;�D5��fS'��"�G��Q�=M>q�zFi[&i̤��wG���w7���RO�T�*�P_��-�-R�|�d J8G;�y�P�ap�}��;�e�Fz��J����H44��=U������ �`'� !]��t�:V�-��Pd�j0�]���tc�2)�Mc����t��(����x�P���@��>��vF2?�0�z�G:}si$&�3�z{x���J�h��	 Ѐ)�Y�߷)���}�
)�NwM�UPZ�R�i-_����~	�dm�VGQk�C�waW�������B~K�uV�=��Z�Ýy��a�sn	8��-��v��(�?fV9d�4�K��wn��	��џ�yk���_��76�Ⱒ:�A�3���ONr��Z
|L��a��`���>�c����jMąƻ�b��+t�U�0=w��yߍ�4�)�n���v(�M���/C��{��#A����W���`Ej�"tZ�f��2�����.����>\P��܏�[�s6x���2_��ͥ/y?}C$Y�3�]M�R�ƙ�����b]�x[���98����`r�*g'{I1�xÆ��!#���G*cETj�H�s�X��^{�ޭou��x�3�dd��:F���Evm��4����������*k��X_>t)��ASW������k��~����\ffe��\�>mOCM���-hZ���B��j�����#��4��RW�03S�q�F�<zT����@�L` �}o�_ j�:�k˂��SIn�g$�>��^�BK_����jU;!/s0���wL��.Qʱ#�o�m�h�#�p���S�������Ƽs�_�ͳKs���xl�V�Q���...��o�#��6%��6��J'lg$��h��v�ŊnN14y�n���v\����K~�l���w
}��衵����߬�Ԑ�ƾ̜�^������b�J���M#T*��GGVƇ���橷pv)���(��3Қ��ٵR�t��R��/�u˺���ݽM�c����jj�em��ܹsQ;cG��^f�մ�܇�p����Co���(�29�4���vٱ�����#��n�LJ�s4�)�z�^�����U�Y���x�h���ԙ��޳Z��Կ?��`��p}������si�Ƒ��/A%����IkO~�-�<�B��j�:�LP�Œu܅	�C(���ޝ�!��.V�u8��٭d��7��s���Բ��4��J���vN��۷�޲���G����~Õ�D�~м�����=�?#�@\RRty��VG׃<�ssL�Ca��l���A{�_C�z+B�D���o���/'Q���wr��ּ*�{>.99fi)+לB��>  ���j���ȍuY��Q��`4K��\�/`d-a�Obbz��J�O*�1Q�Ū/0�l������x�����8�w֙���U~�T���*۫�X[+�{�g�����A*CBC�76�w����܀]�yt�r*BͶ8����{�2��T� ��ɴ���H���@����h�3�eJ�1�]ȡP�g��DRɩ�((-C/�E���%=�Y0a�{E�5;��x�Φj��3Ԯ�H��V�ٝ�F��F�qҰN�����?,�*p7������Z�^�&�sPc'�F�+��p��>'$�$g>���"\��Y���ݴ�������~Y�з8�ˠ-��^ύ���c,}}M�����<;@��~����+���q,e��<ڟ����� ]^+`z�Z�ԅ���g�G�i�<�$B �����\J�U
*7�Kt�d�I�t5�Y���g����]7OWݽ�(z#���4z�`�qQ˷|ٽ���|�Wq7"c��+grJ�l�G�X���T������<�+W���~?m�'�5z���� �#��\�y����w��R�c�V�桡��#��H�O�����S��bu��a"��ח��n�����W�2z^Hf��r�T��!Wt�7���$;�tQ@\�sQ˃���7d���^�@H�H��	#M������'S���e��ގ�_�F��섴v���[[ge�u�0�
��R`��&߼�5Y��_��:a������h�����O�V���R��j,�c4+��1`?>e_����1��ZӪ����9�������Z}0�؎��w�gG�X[[[zxȻT܏���n�Q��/BOWW�a�pCR_-	�������,s�[���P���qQ�#��3mh�W������o�3QSK����+� C_kK�]����s9��8p�Xe�F��hmu�-�܌8���/X��'Puzpy�B�e}�̤s�Y4���6,)W��MP����w}`	@okk����O �������<R>�uvI1r���M/��=8LʎꢧR�h��{	(ϰ*/�n#H�T�Ԏ;�x�����w�DE�ntȿ�LW�<ӫٶ�.�h��Н��_=��B��4���2��V#��՞n�;؞�1���T5B�\
m��Q�ɓ'���=}~V��t�5	�#��]��v')Ů��٤F,�trc%�%ҭ�~\1�tv>ەsY(==�▼^Bj����Uo�؇��?�6�A���"�5�H�Lb��)���:S@ڭR!7f*��h�2}t���y��'ǰ��V,��L�=#�t�� ���-=��4�F}�zn�ϳgϓ���ΏD?Y��(�N!ėC�(!��J���mo�U!��q�T�X�4Ə���Ug8Q�~���M;���� }�K��4��z�Y���ѩ�sD�H�B�����oD1���@�v��KyVS����hv�p��[�e��Nj6���j-��
(2�7d�r,yr�=��B���hԆ>�4풲��8��ړ`��.����.z O��n#��̬/�~�u�N���U�#3Mht����(H z�:0X ���B��-�^�$+ۮ��G���'~Ɉ�������L*�Gt�nI��P`O\0E��ys��}�k!!!��폷n�zJ)9�$��&M�����8�A��!�Gk[���п&��wo�[9w��~�]�y�MΡ[��=f�e���G�����G���_A���Uz&S��塊��z����S3��=\>��-T�s���G�o?�E�=}�4��bc1ף��h[�3��u6I�{��g���d��݇j��x��b�����o����츢�@�_u	������Y��e�(e/*IJ�Ex��CukgD|���0M���%:͉�]c,�#��mU(��gcc+x�R%��ԄGk�|nW��@`n�e�OԨ����ц����V��P���EF^;qQ@���d����lg|�`�#�sO�q��ot;�����b�O�޼����|�5UnM;>�qF�u{Jҟ���I��ƻ���/a�l������Av���hЙ��/G��D,�7)�rA?�@���1z�u_8Q����|�X�ڲ�a�)P��	Եn��5]��Ft��
��b ��HL3#+����#�^��	���c��Z�ǸD��%��_a?�m"�]�h͇VQOR�`��k�3�P�e�*]ũ�$�F�7
D����
ko]������Db�q��LM���F��H'�3S��1> G�9|���&��+��Y�?��_~���l�2z�Y��
���r|&h<����Ay!9��2��ʋ���#����
��ht���Lg�s�V�^�*:�bE�C�j��L DD�c_���,��s���9ϑ�0�ø��oi��G��4qDZ��I�gS7w���[ܾ�z�<q+;{.�Pۓ�a9�r��r����.J�,{���i�Њ@�B��	`�t��Fx��� ��Bd_��<wpV�c���N �O��;�t���D5��uv#S�6��(ѹv���|1L	�={d�z�0(���k�sjK�lq<;�>�D��j��A/d�  RE������D�x�6����ں�?���H��_��ǞB��܄0�(��ȁ���t�ltt� ��v\6^$Z[_x�`r[��_�����ėdyL�=o#� ��Qv��u���7�ޯ�����|(�X�ȉ)Y�&����_1�D��Ց%����'�y$V�5.1ѕPp̕}�d��("����y�)P<||&b5\[:���c̗���1��o�#�-��l^)�xxĉL�d��"N���R&��^���]��[}؎t�X��G��Է�`����H=e��n�/<�ָA�rRQZ��脠�F��� ���GC~�M�ڎ���`j��n��?�E �	��4>���_x�sB���?L��g�\O>7P�/*�
:�K���sn���0�Hol��*a�Nz���0�����	j����W��0��0}��
�rQd�j�P��� 3����V�]�QCm���m�����5�y� �����dp�
�)�ϟ?X�am���Tԁ�xb|����Ik�c��r�-t�t���R��ظm`��%�����C�)F�/������pF�_��� 7�㓩/=��~G4��4k	�Ig}%|t�X6�~�%A�=�;�s�����`�-/&	`�/���-ii����-n޺U���nc*d��uz�8w��kQ^�1uN.�Գu���-�p���d�77_�uo�tء�$H�L��Ҩ�y���3>������ƺ��P�騮j��Ww)S���X�p�o���p��E�P{{����i���C��*��=�SomⰮ�p S��=
��cZ�Mۇ�ŕ���0Py��p���-�|(<Ai�t�f�o����ur.�Ǹ��ݦw%�{$��K��ۮ������<��61{c�>'����oTTL����������b�w�&Q�i�h����/h�R�դM�s6��O���좗&���?O9-_i�by�@��4�H<�Ua���U������X����>��t&�g��6@��D�ĥu��,�c�J��9�K��]1���j��?�E��![}�[I�(��7�}J�m�w��P�����X�9y����S$�>���G�ߡ�A~[�"�)l��7l-k�u��� ��P��w�U������pp�Er��[�. �����\\\m+��Bt��F�ز>�����G^_���OV�_�������0x�@�?�Z�֧ǭ�r�Ŋ�i�tvI5��s݊�T�%0p����vyujzm�-B����L�ׂ�j �er����#@x��~��.j�@(��^���������g���vg��w�WM�A�}#����v/e3+�1�Z����wR*��
7ޖ��zz�@�x�nG��Ok'k�lA-B����M��>q������VC�����~B��L
7=~Պ(}��J�*�!1Ҋ�X\Ӣb������bX@��2~u}y�8�|�{ѹV�u���J����XG*��k��Fj�ZaT�������mċ�_�n!��/��%��zH��k�A�1fbh8N��=<��b�^��_
[ppp�yCX���\a&�(���׽�����$v���߮��k�+~�V���K��Y����XZA� �?`���Z�5�s�������wɊ����]��������{�õ��Q5>3}`�.%W��x�!���ah��ŧ��\T{�*�}���$�%^�0љ��K�2pŐ��<3N,��O�c�s��'�g���S-TN��肬�ᕠ�w4��� |���M,O����)�Gl�*ޮWbR��m��Q'���0����W6���^g��P�A�ر�sjk������Q_��Ovt?�ʣ���O��F����q[5��V�5wC�!��%��Zj��ړ��n��a�0����"��	ﾲ�2�z!<.V��qQ큚��yi^Ŋ���Q~5n<`�0h�����L
e���-u�����s[Cö�C�g]���(��"'�nˍj�i8oed�$m8f�j�K��@��>�Vy^��qdE���8>� A�@X��In�`W�ĉ�9��ų��A������.#A#p�}۶o�90�_��Ý��({F�0�9�R�t�'~Gw�W��C6�����AIi �yD��]���"�.�̶I�K	���[�������l��݃�XV�Rv+��&^M��3K|�p�V`���t�����8��h"�~b_PF�o�k׾ж�ܰ*�$�`�{�+D]YRv�K;��n���2�	�����(A�A+noG�pОm�L���G1�c������6颫$7R
w�������Z��=��2�"E���bԉ�73H��wڞ�G�@?f�=�yAs��?n�k�!�>���h�ހ�X�8����max��kr]ϲH��B;��%wG����l�&4�������%��}i��=�A�+�4QDih��-�1Xf�0��~0æ��)lR��;~�x�F,'H;���y���X1Z��ʅ9Wd������m����ce��un�^��i3�c��>�&��E��{��°����b�3N�<}������1>�k�Z`��\�]�^:[ƾ��%J=��ú�R�N2��}ى `t5�"�l�n z�Oa�xm"i�M>zs�c�	�:�1��C�)�o!�.�[�p*Wg�L�L����rs��~3HZ��my���]->>=���0{
ɋ�����<YɸP�'�}@^����U�jC^�y�r��P �����wf5��9߇+
�K,� �K�l[5�)?M�PĻ�٥��+��y���	lа9����2��9��F8���SfT��aO�o��0����M��"��E7�&R�+� �s��ǹ�1�Te�wnt�Ӈ�HF#��o�;�Hq
`�R���|����̉�s]&��g��T�t�j-�2����d�I����:R8L'zJS�B��q�#^e/���DgN}:�R%I�:�۟�{��c��?
I'�ʦ�3o3&��o1�o�u��sͼ���2��m��t�s/az+������}͹� �ii衙ϼ�e����/�*�x�:8Z˯nNB��U>dd��j��՟G�ج��n�x$%�K�&~6kg���_� �uݏ�����lEP�7�\��N� 4�ҙA�"
	���6�3q\w�m�=!�qκ4L��f�ƚ�s�W�a�h�@��T���f��v�4��n)�;ww���YI��)�|�����ҭ�֛_ �Oc�Q]�n&3�տU>+,��3n�	ޡ��B�k���T1Y�	�W�pG睵j�� ޥ�9}�Ѽ<<q� ��{��W���8`�An���@v�6�\��i�c�z'�.J[��fX��	H�A|o��Z��y��s�eԋU}��E%>��DbU���D����[�#H!�S5;�>���|���c�`��Ũ���D6�1s+����Wȭ� ����E��q�:��r�u{�^\Q�HgMy����󝬰�v�.$Ӟ��"x���%57����g6˝�<���Xa�*
7:�qfo�7�%�?o<,�����zf���I��},������^vY9V��	�(|ͭ��"JPE|�!Ӏyl�2���gC�S��]��T�n �����R��Q��S��nHd.Wx7�gʴ����릔�����!K�u�T���i�ܯ�X9L�@v"��V��K5,mЌQ"��1�x&�%s����wJ�n$(�
/TUn��PhGv�Q��OwD��?���#2д�h-Ɗ��t	�a�N�����_�hk��\>�Т	0{����g\��(!>�WD���@a�j�֕����c=e0Pb���3n���a��7���D��E��Q���|l�J��Ġ��u5���L*~�:�8��~�����3�Q^WO������5�@D~u���yp��Ci�۠Bt���Z��{�0ۆ֧l���Gz�~%����i�� 8H��H�#��~�^|�z����@��J�dk-��k�����)F�M�C�4�}%7��+���L~@�
�w+���$��{�	�~��b-G.hm/@�Y�����;>�k�i��nA,'%-�K(L~���S�j;�4��.���!xf�O��3.����C܈�����K�ԪydV��tݪ]��E��� nT���	6�T�Ǯ���St.x|����k����ۄYr��r���Z�x�O�KK;����Z�=U��!��>o�5��B ����69�&F}i�d0_��VM�pA\?��M�)�xORC�b���:4�dt�A�;�q�(�Lg���G��j�u}���
���5���9%Co�ْ'9fQ=`\��ߑ貕�Bx�4���>V��X�^
����xW� ;$f���'�T�k@:zw�$�����w���n����2��/�QJ��0�`�lШ_��K3�ɕ^�����KS?�L^2Q���:�i/��O�	nz'~��#������g��+�IX+S�`���/��},g�Y�����_a��F�6���]o�T0��c?�L«�z�8��zh��gne���7V��*�遜�M�Q�yc�5�'jo��6�)S<H�fD������_c��4�=�-6l4/^�R�s͍Yr�6�:���T��O���ؕ~E���H�6��N��8g^���T^�յ�z�13}�����1�A�N����p�Z�[���q�w���"6�̮����L^��Κ�<�`A2Ȉ��� �K���d�;drD?�Zz٩r�x^R����B���.']
)�������2��'&��~��Yg]@$��Uwd��n�03n��v􉶓9�W��1�����#Ji�]]]{v�9��W���7O9�L-�̪A�V�EX�\�;�:���_���lgg����MF{�0>o�Kωu�R�h��ұ��;X���СC~��8�:�}5r����s���6�O`fS�N..�W
�cX�5 XrL#�����x��XN���p~�U5g�<#*�W�ֵ�?���Z��].���P��P�������3k-vXQ�:�w0KVFf �i�].U���<�`�9,��}��կ�Æ��oq�,�V��Rҟ̏�Tę�1��{�n�:��y/�7�&^��t�������.��2US��X ���.`�ծ,���+@;1G;i�͑hu�ʂ�PԈ�o͐Gɮ���v���$�M�-��>@���4��@�<P�G?9�yk�)B�^��$�;���{3���[RR����a{{��6j� ��_��6n��5�+�-9N]���&����%O�l��J27��od��ӧ��HZ�r?��	l��m>9s�g���e!�I/�#N�{�m����̺�@X�Dk��7o����a '������=�����Q(	�RD�y�ͺ>Wr3����<jq$9�n����SR"2a�Iz���3�_v-�`'U_��o�ju�K��he']2�^����γVb����N�ioI��&��\�o�:�_Q-K���5�r{aҏ�9�5�v�ơ55��3�Y�V7	���3���ۚ���y�@P����|3��
�ؚ�Ȉ;���i7V�����\ju\���]�r���m��!�9��=�$m���K����ls�f��'b�(Yy~olM"&����E��.YKٚgIJ>�7{��dq�x#/�������}���F#�����m�zc�ן���<���A����|�ԍ�F�k|^�p�om�V��Y��Ɔ>���!L�JNd�u`t4Su3��*���qz�� D��y�j������8l�������{э��0sT�K�D[>`4Z��m�Sئ���K�b�f�L�����K�E�����9N��&�c�s��(�^���2����$g��P�4��H�kV���G�NaI�,����/~+��U}�<��+��µE 1<c���ߝ~A��[p$ٸT�8p0~ZC��ew�V)�FB��o��t�  ^���A�.d�S_��8�Ҝ���-�����vϟV�+Dtl����XI�Z�Q�<��q��҅��ݎ�'��H#�& "}�=�9͎��y����j����@�e��@q[>�b�{Ĳ(�
������6�K����H�?.������M xB��q�ѓ"#1���T})����t\U4srsŻ���u2@��
��v���nf�jr$]*�|��oڹ��o+6JWbo��G��xV�Nk�� n�H�%����5��V�S�MNճ>y�D�)0���ř �{��]\\|M�m�@_;tSV��9�#���|�W��r�Q��^=��^}�2cԔZ�_��MP/}�d�g�넔fh��I�8:�_��3���/9n�Sui�n������F��O���^�*)qD�Y�D������㕌�R26���$g'��H���'�#�~}z~��������e򿈈��JKJ|��u�H�u�~u^���H���6\02��)����T��n�[�!$2�8��겚�k�
�=��7�.[��Ġ�h���h�A�r�e��=�x���I�/B�9��%=�[�wMїsvǍ��z����C�;8W&�@9�Q�ji�������~�(}%��g�k�P2�pƝ�����n�a�5.����ʂ��YD��Z�_��,�@�{1�Y����K~Р�:��Fo��)��':�&�g����)������u%n�_"Z����t�GS�'*�9�0�4o�-��5(��ϋ��Tz�͈��{���J�(�Yj�.�$Ž�_��4�4kd��&0R�pj���1z��Qa�����`,�q)J߻)6v̙���j��H�����&��S�X�T���ߏ��XԄ��[]ȹ?�,�����;����s��C��$5�ǩ{���^K�������/��ء$*#�)-++ہ�K�2�@� ��Q�!7��xV>���-$Q*%�-R5;�C)Y��zbae0
�}�`)��ۯ�
�Ǐ�2��{����r���Lė���X}��oAB	J���9��[�Xc=3�b��\C�<֊lJɪ��DkV���U���-�+F�)����yx����� ��	�KO����,_y�'DPz�B�'�ka�9(9wDaҶ��ާs�`�5����h`��Hp�zK�vy�:z��'�B���_fI��1BH_�~S�s#�A,�����*_-����}ɹVܥذ�}��g�n;����b.�<I�^f;���+�z�CTSH�{S����ߴ(�,������C�3l�M��U0Ӣ8�XU���2��%n�;�ʱ�����  {�"��}]�2c8�o�^�֯"�wu>_<�b��j��7��(�|���4<�ф%a�sw��J�Y�b����Q�&�KjE�Z���j��봜�Ɯ���V��B偘��7����ʮl%V(�<<S�����fF�KVv���V�T�Ұ��[)3#���+-�>[�ib�^Y��&�LI�`x������eRyAA��?y1+}N{)�^��:r8D�[rgg�f�>;�qb@ro���dRZ��yx��ʟUC(��+�̤)Ig�=����ة�k����qXM�8ݎ9��r�d��!�b��}B.t���:�t��{�[��}T/����'���!�q`�eCT��޽{�m�sl����K�<�a=Yǽ�����\&]�f���\�#_�C.�n9�Wb�|��K��@�/P]O%�D]�|��T��+��𜝏�ȻͦT^!&sC��w�:��r&�����L;^+���Q�㏼D�af�(B:�%�4�|�5�W~L��2���~|�<����<L.����Kt�kӨ������@�;�N3�x�a��VG�r�ZWW�aZ�Bl�S��r,?�J�і�� ߝ������W[!�Q���2A�@E����v��C� ���nK����)��+��UA�-Q"�hʟ��i9�j<?��P��r�c~&��)X�>�mb�+y1-�uy�G�2���?�N~'���e	�yG�,i`- (g(����FL�v���ըC-^bFV���C�}�Qa�|�^�!TA37d�i���]�*�;�x��5��Kr>��st�ԫ$N�sIMʴ�Ӭ��u��ϭ�6X�s�u���8�����(�g��c<+��8��9:�z�m�.�kb'm�صp�t���Ȉ�n�D;�׷O�F�=��Zk񲡻�֚*P'+i���Ǘ�+&K����j.:Լ�R��Y��f�Fϔ���F���r|kW����C�(}_tb�n�^��� ��*�V�Xi�u��)��@�q�M��O�m�����P�C?���q�� *�����)�� k�;n��p��!�*���VҐ�FzR=̪��`�2����f��7z����Ml�5�i(�6社�s@G"��W淾�`���ذ/�ᚗ�^"F{�O����P�� 2��tM'�J9Č��vs#0�{�q�<�k��i|?v	��PMO�?�Zp��&�Ss��.�ڗ��j\�a#!�~�ᆫM��Ǡ'{�� `�`��Bj�����>R��$'� 6<z��hW}}}�[$T�ؿ�%���.\�*T����J��]ϗ/���eW��j�E3^���]J�`o|YV�x3�IKK�r�#��֯��3�uW�̖�Z�A�n@$	�IhI{�^�tV�R�y�����ݡk."#�(隽%J�[�l{�އ�\�4^�ٞ�����|�Fn�����$'���0b��ŧn|_��T�
W}׿B���N��7��Llj���Іt�A-VB��}ԠO_J��*�3=���.kU�����[��yՌ;u�p]d4>_�V��5��`O�v� `Cqׂ%toÖG�s:��I��@��
�w��ڧǽ����H'f�����'r�;�;�4J�7e4�)��yR^��?タymn��'���p/��U�2rOU�9냩��J���K�"gZ�WYQ�-�6�W�}|��Į0R ��f̴q&wCR����ѣ7�!��h(}��+����Ul4��{��E? `M압�Q������ڢ�.�������'����i���L~��lx$p� VUl�Q{��P1\͈J�+�pW��o� *i��/ۃ�l�>���.q�X�Z�TF:��^�ȼGe���<w���q���ku'��z���]B��M�ʡ%�\������8�kyz���3�D)`H����6@����23���.cͅ��vX+��i� '�qw�L���!��z�!]s�BS%LO�&�!�a��v�}��̊��ZN�k׾V�׭^��ϣ��M�
��h��9��?�z�ҋ�ڭϭ����nGb���~�d�Jh�0I�rD-�~&X��MoWVF�WFT]G��$�SOSS�s�"L�a����9�G�� h�#v���m,��:���$�!�9/^��?�N��j�Ǡ���]i��'6����q�h8YG?5 _m�¸��>�_YD�s�qh��|�=]Ϩ��!�Y�b!�����{��88L�ϐ`�.k@{d� [�ێ��޽��\p���gDFnC��{�v��$}��KzW�gX@b��<ƒ�އ�싻�����u�:\�H��KƾK��T|:�BN@���:��y�t-�1�\,�����`	Yd+��=ܓn�H�U7��1�����p���<Z�lF5m�^�k�D�̑��Gd4Vi@�F�}_���0skX�5�%?�g+:��DV��'�J� �!��f��Z�r���Nϴq��7���X@�z.C#0�̏��H�����E�r�91I~:�[��?z��x�v��:�
Up�)Y����`r^+Z�w���O�s�7����S�f�N����)�ރ<�)�%#j��h�������AC�ЇҪ\�'ˁ�H���߁��`�O�1��W����C��%N·f��UzP�ǿ@��P�墓�{_��\o�?Wp;hVI�����Hn�/�T/))AG:I1�_�nU�M���B5ڠ�hL(�]'>�'wu��1�A���^�0���u�!o�8��S�ndd�v��	�]�������-5o9�&S.Hvt��u�(��t_:��vh�H�K�9=��۠
W;�����,>9��n~q��jm/R;�&tU��Y{e���Zs߻�Y�yu�q��VUb&�9r�"�h=�k���+A��.W��B.���"p�j}�}�_�i�>�8p��sjI3�.h�o��te>�?/��N'8!�ov�f����ʸc�9u�֞����6�\�[��?�]�Dñwa��ݚ�yϫX�S���e��7op{���w������r��Q���7oޜ&\�mv��Ә?j#�B�_-�{_>'�*"�����������Tty�DI�(�x��ɚ aM񋐌���>��ϸ���\;e�Y�1#�/l�:S�5F;����^X^H$����?3�#���s}�P2:�J*��ζ��6�D��ڳ��&#j�垿W0�Y�����.!�����~ן����v<cd�K[D�)P���v(���c���,����(v�'�Z��
�Y=D��c?��ͺ=b�Β.Գn�	6�{H�BK�Pd�h9� m�5Y4ck!/vp"5�L�Z�p�#	�@�nAГ.󔎟YD�ZIE�����K'|;�#���f:B�wF���z��쬄f� ����B�D���1��zM�vL�6g0��r[�����0���	,%�6�:��+���~�^'����ַ��y�Ol���w�"������V�v3�D����S'�����999���g�mb�z}tb����c%+���"_��%�e����-�yé-�\A���j
~y@BV<+e?K�:�>��]16�݋_މ��ҏ���UX��m�iZ@[��`���%���%%�GC�A��N�j����]<�[�L�.��~�׀P:��F�x_S�֢#�P��$�F����I7�[؉���kRn��T ]K��B�0��)��Ϣ_��~�W�&#+[}#�x���W7����ܜ�㇡ [ ?ֶ9��%�ݷ��[ODT��Je�H������7á�s�%V����E��K=�j*�g�5	ߜ
��)�����S9��񥠷��1|��p�����En��(����l	�硟�F��o�O�N��~7}�&yA@�3^�����4�郞P��p��Y9�GzzP���+.~���}����nk�W_�N��?B��;���߂�j>G�W�Cy�̟�_���d-uX1��`��{\��c�Ⱥ?/��g!�|G:	�it����x�jq':��twÜ�L
k=oߞ. ����R��m=Z6�`w W8$��믥�(?��$��?���9Pp���H�����Ë?�$�+�nz�4o'����6hl[��itRˉV��0��̏�ƐY>���
-�N��+�d ++�Ld�s9}�tr����g��j?~�H�ƅ@z>g�v��u7V��(R��3ɲ��Yi$)L/��E�eu���B��'7�J���ݾ
0�]�k,$)O���8�v>�f�w��6a*2�f��t]���V"�	3�j������WǍU'Z�<�]���w�c��ٮ��5dP����P���f�z#�]���y������%�0�n�7b�_��+��U�6*:�/��i�f���O�A�������"\�Z�ZI6]�������f��~E
9/����(��+n�*w� �.Xh�DA�w0�{���������k�BQ����[���w�.޳{+���j��<Ǟ�W;t���)��]�#���	�X������W�It����`��YOC�(���#TI�?��;������3*���q��b$�`D�
R,�:D%*��P�m�Q z���Hs�л�J���;�����?�g09��}�^{�s��y����0��R��.���C�:F���ky,���������|ӫ�7l���,�����j#���8��������}J`!� ��n�$�j���״2)�d��-������6����B(��^\��ҵ&(��Tjj�M�;� �4 £ҕ�c���>�{��F;��(P�]�����VƦ�1�Abo�>�R7���cUzi�b������9�)DB�lQ_��H%�F��vU;�؅?��c�ޑid5|�ԑ��^ �U��DD��9G���UxJ=K�LG�`����x3W�L]/��$.]1��	õY��\��'��#F0�W�2[����p7��ύ~�*��K,U2}�����f��X�2���=Dz@&��<��~u�+X�/�X��í�?ݏi�K`��B�NrC?�@����"lM��o#����HD��#�������^���u}�k�\�����U,������qo
�ajS�𠻰���Ti$�"�f<�a�:��@e:v2|�3�;Us��~MSǪP6��4|�)/��A+sC�r��ז.X~ìO��y�s��������:X�Gw�ݸ�gJ��߲�v�A�!���]\$X�ښL���^\��������V�ӳW�nmc�]G�dcx�V��qǐt����"��r�)�{����~���*��5��D���]E�WݣY�n!���Q�W-�M������W��pa0�SS���;`zƟ��2�o��ߑV��W�z�a���T�4��Y�T�<�#e#'��*w���"�տ��0,�������M�>�)�ǋi�88�ﮘX����M��M�R �"m!=B�B鯖HJJ��vbo�������3�F\9]�1�뵫�M��(b���/� �7����w
< d�.;�=n�C=O"�-0�O�>}��ԩ�=d�-˔V(T�=(�"\s��Ks���Ay155ݷ�$���gμr[��ҥIKό ���c�u)))V|��b��S@���~�$�Y�Q	A�zf�ŵ�o���*Ў.�D/�?�8$*���,)E|�
�J�N�j�8��ޠ�"�%j�o����ɀ2�crL�����P��W��\	�>	�s��b(���F��u��n�惂����o�cg'���@������R�377Ov��ɪH���}}��N�XD��?MN�r���-�z�������i��Sc�^(	.�[��@��I^ЀUJ��h����O�� i�~�wr>h1	�%+���+����y%���ϑxԝ�����[�`:�DB9��+ 
�Z�Y
���gd|Ϝ��V�<�нQ�Bi��ڃ��7���y+��.M����*����J��@7�>c�&�[{Ztq��?u��������Ҳ��vHW6����廒LW7w%e����R��n�tO�����`��C`�9.Ns?��H�l�"i��>�N����)C+�O����'��p�e��_��*GRx3�LPV�}��Ý0�1����
�s��� �����dg��ݩ���^�Cȯ���6l�I�;c�+��lI���*a=�N����J&&���]���~�p��!�z|k۝�c̕CX�L�^�U�g���ݲ
���xiD��Y1Z�330S]X�2��Q��C 9����lI��$#a%k *�c�)G��Pk���X%����=��=�$���T,@�.ɩ<A�c
���Yg�N'�|�u�i�r�#Rʀz>�17��y��n���!�qgT�ȄZ2�t7#q��{���qRx���-�/*?ӥʣ�	���9X�6qRH��tP�;�0�<h7n/����-�
�G���	'�	9�p�P��Jj�W>�xz=W.�tED,H��Y�q�b��}����b�P�i�A4��hP��)T �p�����b5.~[d��'*ߙ�� �^�-uv1\��A8��W�5o�ׂ���m��w�K>��z�ξ��*q� �mu+�����?�-N+�����t"5��=�/��իI��#\\]e��O-#s[�G���[�#rW�}T����{fN9�<���A�Ǧ�A��CQ3�֯�9Ԕ��k}6?feo/H���p�W�_�Fqt�fD��2�mԥ-MP 22k��A��6���"+�U��E��Q~������-��+SYiu�4���p�`:.�h(G�P:�	�LA�,��K��}�Ľ�����~w#���"MtoP.�ך�A���e�������swR�r�&VcS�ͅ��D��o�J��UP+a�,�X��2(���oܯ
�an��;=�h�(��t�)�g����H�d�SיA.�G��B���Y}dsp�3���%y�Pڃ�1ꀥ�� �p��!ٷ�K�� ��``�Q�bf=�2Ҕx���=�s1���T�.�@Մ2�%�,�x�QX�B�~	?z�J\�k_<Ճ[��(��[L�[��F�aѭsHˈ�sP\5��ǜz�p21ȡ��9A�b��t0w�ӳ�C�Df�E_g��c��k�!��E�E�KVR(��#sT��qJ�&���؈�׷��ݭV`e΀�;���N��"�yx���_��\q���gE�B����RЮS���@Xk!����P��;��+?ruq	�Qq��(�Mp��
3�+6j�#�(L��y��́��Nl*�^�?ѿ QΗ�M�v'�Հ��;/b˄?]��Ugg�]�N-<��z`~�԰P#�0��6�:_�)�Q�~�������PYJ��V��ҢV⤶H` y�[L�4�Gb|V�튟�Ӆn������Q�n禉����حx�9�L�s[�\dPQ�" 4JEK&rm!o��%<������-_?|��<տʠ�U��'�k��D�i��`�@qa��͟�i�œ�|M2V�P��/_�y�HF��������V&J�֚͛��MO|t;�#�D����#Em��+��]8��>pu�z����YD�Z�B���AF�q?ݒ�ϫ5�4��$��`rې�6ʲ�������]��E��p��l>��9uK!�Y���nNؾ�DDF.��\�(��t���1��Y��>J7�j*�`O�qxOq���2�S��sH�t#���Ur3X�;H� M�����
�!:o!��zᎺ(��	��'��׽��e�Ց���+A�?�,�YL!>��E��Q���[�f����XƁl=乸0?�!��["L����9��
nU ډ��a�/]�7Q����<��#B�ŝT��ݭ@�aK�/1v��sBQT*�B����q��lE?�F677w��_�o!�$m�bR��l�����q�Peb��~���G�Sp����l%.u]�L��xV/���2�{va���Bw&�9���-�\�H3�W�\������j��r��rBI���}�s�a��`�Iz��b �'���u��x�>Q���Ah=
����~�/OED��mp%��B�b����� �ٜ l�Y�d��+��zq�ዎ<��i�F���#�J�/eD�<��u0���2�'�!�@�^������c�ߑ������@��� D����Gc�q2�ᇴ�R��f���>4X����H�
�L����84�xҭz5��/$Ǣ7{�Om?��7r���;���8��w�D�{<��a�����	��W!���G+3��H���wK��RV�1I�ktD�97b�b@s�]_�G���Q����Ã̺��j�F�P��BZE�7*W=�B�Ǭ)N�?@���}��?�)�MΝ�Y�J���8R#^@L~V�v��-��B@�I`�" z]X���m䠯���ᑴ-v~�i'qZ�K�a̡6~'�
��)u�3থ�H0a���������ƻ����N��ܿY�=����`SŲ`�6�`Sf�$i�@�L��{;c�̙ˎl���{�9+����?S4��]jb�y�:�ٯLԞ/���F�+�������b̽��Z�\��v��}��ǐUiK�A0l�/�����b�޺�#� <��HI�D�'��� ��@#��oذ!��O|BD�.��X��!��ax���ҫe�k��NT�ĳ�-�k����TD�2~��b�45�C'84��H�j�koޟ�M�ɾ���Q3��R��k��P�
�;w��"y��K� �y3�f8.}m?Z?���R:8t�)�b����ԩ���;帀WpS$4p@����Q$�zH�D�HPg���lGՔ���L�Up�9��߼��)o�53[Yh�9p����#*�þ��x�*n��x�������[A����Zg2��F�[��Z�WX�Ȁ�;N�LTS����S������n�'.fgAʩ�/��B����Fr���ғY�c�O��\�~����@��V��@�5Z�P_lf_f������"��>�s4�����,��b��\/��讞��7��/3RP8xA��'��͗�o���.E�ϻU���H�ə��[�j�6��*Q�įAߟm�u�*]>H|�L+��j[��3\z��z_�u)
���	|�o�mb�s��XM�D�W�E �o�+kL�EjQ�� �lg��DB�8�ĥɍ���W��[�8������w�|�<H����-A��/ޟ����f��}�^�j�S)�Y(Ҟ,����I��2����:���:�#���<���4l{
�Z6g�ե��F��4���9Ků��S�Ʋ�7�y�*{/xYz3%���d�v�\ڶ'�.�%��L���>�W�?�o���"���q��('�R��R����:i�Ny�ˑ�X�JH�\y�~	�ҔC����,�o~O�͛�e��d*\�#E;w�:��C���l�z�0�E��Yr��G?���s/�����ٗ��J&��Vimi�Nw*ؚ'`�I�q�z��fNyC�W�|��k�Xzۀ.0ǚ��D:t�P[�W�Vi�E���̝W��)B���r��tK΁8��
��Q#��>��N$��2;?����g�>�wV�Hv~$y�B��]sL�5+W��bs
��e�,����d~���y��n�}��9`G�O�����Qv�dXeE8C����9Yخ#C9���+�B{k���ve�4����H���:W�ƖmR��v"D��|� ��N~T�|VW���>����k<���" ڟual��`���K���Io~���_AE�Jy���&v(N�6��}� �nla��g!�9��<΢�jK���65���W��B�9��.7L�`N���xБ����f�z�4I�V=$͵�d�nٲe0�� V��8Ln��.�Q�x!����@v� -'�j�^^I��HM�Ӭυ�A�X��V�@�差_�fy�}��	�����4���B<
���Y�6��V�©��퐋���"f����Iĳ�ɝRi�ă�����r+�:�BCj�z� ������ۙ��:]�.�v��k�e߹
�G��=x�Ţ����������hH�^�r���NYM�)P��jjj�n0���06ȁ5�_pdO	V;~������k�l0�&C�T+�wD���Ź�s% ��3�M��Y��ѕX��q��q<k,M����S#����W<�H��
���899�:���V���=U��-F4�a�Y{�SJ�ɰ��d�(��т��10a�H�G C�����t�����y#��"Iu��vJ��יu�%~�R�>�������1�G����-�⣋��>��-��H���oϓdג�@=I�	_�t���c����dW�'�P�-f0��эFFF�o_Y[�	�{��	��W����o�&�Fn�:J~k���H3���� &&����R������z|��OTTT�����x��iJ�o�ߪ<������q�9'��w�5L��=��^�4ʣ
H�-B����� ��(x�l�Pd�*-Z��'�8 �r��k�q{�����ǂ�u�=m������lF-�ug�?���c�P���{�!�s�ls������΅�~F�%rKxIz��2���6Ah��ܽ{7�h\@I{+j��y���(L^Ԉ�����=�9�!Y�"��)(k�OTtڮ�^e�)�j(�<��j��g�� �(�>�Xg��������ϯ���y�Ef'�a��=UB#6�nejC�z7�xw5�U�Ԓ[Ԓ�\³_!xC�F �U�sWQK�c�''8�w��� z,��ݻz�p�GORQ"�΀��~�MO�
�ȸͪb���7�GH!I������i��H��˅_y�-oy��ŋ��'�}��(�Y}�����+p� �%��&��/���"҈R��ACVFƧ�0�k8_.���ԝx�@س��@��SVV�-.����p�z����%���9F�ra~�H���)�J�/�U�ǏȖ$N�����SE��mXG��:�sZ����>on���Qp����T� �`�o�cb4)�|�f5Qw8T,�3�N������7W53;{��VVtK��@����Ç�]'[���l:�$�E~��`��~�t�20~2��� dIz�Y��*�w@�Uz%rXU,�皮^�:���aD��8�ڔL�U�q�ι��**+@�?�D��-Y�e$����ŝ��X�ɭ�C@�� B����;a0����c��¢/T�Z���{��{(Q�8<�����>����S�u�n-�[��;|xD��L��m��960h������f}��Z]6�s�H�ZZj)��~!o~6k?J�_`�oB袓y�^?:kTI�������&$$�F
qe�Ls�^]�(���R
�˼��p��;lJ�F�ts�%���탨v�ƞL#�Pu@���Sq)@�u�QXױ���+{	ն
�&�;�gp����JX�d��jn�8��W�\er���C��gv �KG\ߣ9R����fef�g@~f֍��ui��|�(�q�R?uE�p������P�+I� G���e��?�u�+^�vS�Z3�f��EGvk��J3ss�u�W6s�?�I��a�]A��9�D<���{�QX�n���_�par��<a�S���؈�
J�Y6"ۺ]Լ�Z�b(HzU��{4WX�N�j	w����b���$s���1	���̤�Rc������>��kI���¿��N�i-7����jr"�]SOoo���c�Ќ��4��A.D>�2��+k�2Q�����W��W\]��^l�pΔ�j���m�B�*�H�r[|s>db":5�y5p�q�)l�H6F�w�&������?K,������vbJ[Z�Y���k/�/A7�r��7�ڜ�����H�����ȝ��34��s��d��Yii���N���V��<��迁��v�'��?t�8�#!�3�M�J\􃃅��5��wC�[[a:Lօ4R���]�v�v���fسP��k��L��A�Uk�Xx�I��D��ߑQcH�
<e�4��i�N!�z���~<�c�#lX�b�L'�����{���x���J���ѳ��+�S-�d+�xeK��,2�9��N��6o�s�
����_+�p��������4R�[���ڷg��95{f��\r��N
�<\��?z(ܶ={���z/����q��azO�n�h]V���6�P777�?5���GVn�̔�~x�ɨ��x�[#���B��Ke`��wp�����C)�%��Z#����N %�3��~m�ǉ^��)��eo���4�^zr��=e|��5��|�̠�FJ,�]�"�C5���}�5�5K0b��)6^� ��<��;(��7��ٙQ]����jei����m�sPw)K��É�7����QS�l�'q"���xfI5M���������o�)�E�`XeX�0H)�~�шς��;e�e(�f�f��=j�Z��o �wv)*j+��,�yL�v2��u�=j��4
C��7�*CҎ���U����w=OJ�;�3�GCB
g���}�˪i���ϵ��4��ݓ�	��U�}�|M�B�K�"��I�A���,1n&��KSs�_� �D��so�M@�CUcd��ۣ��Z�Kh���,Z�Y�`ӹ/�q
5�D^���IYf�W�VU�ă���r�w%%%bԒK��3����a@�h�Z7/4�?dn���4���/�^�-Z�8�i+��~aFU��/Q������s�1�M �����pH5��)	'%%%14l�. �/tB��~ # �W"�P.(�(-�ZWo�%Z|��a�cPѢ�#ۭ0�������ΟE���[%D�{�RtvJ���-B{��}�����s&N�lR��f���Vj#�	@�
�fJt�_��^b�������f����YR���5t�Dx��RT(_Sab0͆"�G)Z),�!܌c�?=[o�[x^�u���9G����.�����ɇ�_�\�3����2��Ȩ��#��v*��h�0켬�c�5����i>��2r���������O~<ofW���}�{���;w�.y�!/ό�p�����>Q8Fr���x�|$\�|S��qJα� �� ;�U뭕��Y���Jy�_��Z&��[?ۀ��!man�o�m��`���tFx�c���l1L��_'�O|�	��iד�&�}pҗ@�*��@���KA�xG��ߔ4r(yG�^�U�tyB�5.7Vkfe�>�oE-��������"<}�c��&�Xli�낧7�[���2)�@���Osdg�}e�ы���4`)EZ��o����8?Yt�̙3&�T��1�vM�g�X��5[�ju�zw�(�xFE�%��Ve@9b����z�/�0��5�4WOF>����ҁE�%�VV51;O�
��B�޺�ufVP�3^�L�7���_��whRL��V�jx>E�EX�#Ti)�*��;��N�LKm�T�p>$�%��C<++ַ�>�SL��P�b>����گ\��!�.�[�*�k�+���Cp���dKMɰV̸�hW����
o*��ܙS��!����ВZ�X��7?nK�G�Lbxl����F�����ʬ|gf�(A&w��������'��h��=�[z��<��)|��ķ39o0�:�wԍ��/�V�ރ��-ya�{��9��+k�}����F"!#��̬<�=K,l��3�+H'���Ƃ�2��ԅOh��u	#�{y+��I�s^d����p��
�z�>�!��������)�S�sG��>�#:_ݙ��=�n�@��S�O��.��w��.1�H}B���K���dwi�t�G=���R�=�2��ߣ�Y�:�%�I�rG��ϩ@�����n���
�?_��i����x�-^�沦��H{�����H��@����C!g�ܣU*���-���#FFE{�]��7����{@��.)t;`���+LB������-�WW
_�T$w@����/![�l)�&�|h�-�5����X���@ԋ���ڿd�׽�LI�I��$���>bae����a� ��w��2<|^c���/�"�oOe��6�y �-|�[�tch��S9s�?}biW�O-nPڭ��K�ܰ<T���EmE��A
p㊞���������=fS��\�5��͛�WVVN��z�(�+iDo;� �H:�$��^ā{������`V� ��`9�I6� a��:yN��K�jZ4��zlٲ�R��ij�cTԶxqDr�����7�.{���U���s�c�˨��sl 7.rw�S�x�:��8�O)<;n�<W�U����7z���(��Y*m�ӑ�f�F��i�&������\L��n��)�*�,�E�^�����&'�F`��_�::~�ĳ�,s�--AR�$��t6��� �X&��U��&���A�pHc��V<n�:tg�Lf�CF텀C*;�8�G��"��0��~M|�P	��v/�2{�9���G�S����)��}�;����NL�����΍���k���� ��9��ݷs�ab�y�
YVC����#���ꞟ�J�g�ey�
��y+t�g��h|/
���&����v�?�k999� ��X��V-g�͞��t�$�p�.BX=g���4R[-|E"�o�7�?���/�)7p����( ��4)g������� |@<��P���aNu�K���C!\�i�8���c��Ω_�N�XGj����߿';��J<R�eeY����y��hİ&��o�tD�E�@~�2��`Q���a+��<��1NNIY4��r#A���L��@9���Ņ{�Es}�J���9pOMm�x�$��$f)� o��U��dT����"������.Ϩ��}�D+�7�s��,�㩌����F m�SU�~��{�.��|��,��dl ��0�6J�1�B����O"��h�.�p
�,'!!a7���1�E���U��a1��㩙���D(9�ImCVp{�b�9��`��* ��U��!����۠��x)�-s8 �{<k�+��B��̢�9��ҫܞ踸��L|�g�tȯK�Q'���G���A�Y^'�����Mg������^���s���K4v�uh�>(��q�;?�{��P��.k B��L��*���~�u7�<C�}2ӹT��,Iz��ƨ��
�#�C
)���e���m�0O)�����5j�v9�LAV���9/=�mR��

*��_Ak�#�(�HIe,��*�(}�4�zʠ�!�a���%���d	��(>a������R�HX�SS���PRU�%̺"h�D�f���'�o�6�w�QƘ��0!�N�(O� �< �g虝:U�`�ߌ#{\���N�%�,�"��r/�@�R�h�`�|�{2�X��c,XS�t�s�-.DO�;�'s|I���R� tܣ�̂
 �~��N,�4� ���n<6Ч��
XCh��JRҊ����U#�rR����JBB�	�R����d��J/���������>9���O��**��Kn��g����h�~d���3����)!�	� ��f��T<�鐂"�mR`Z���o��EUYY��nI:L�����0Yqa�$����d.��j%q��Ϟ��T�fNX?E �@��9�Ü��[���d�W�iDR4$eE�.q�_0*�@α� �#S����A(,�Y`b,7���������W��=��	cc��(��(^n�w�N�,�d��R�Jͱro(hΙ��%r�S@3��\�R7��r<��!�I�Y̸�� ޓ&�ǣ����
9g'��ե[�IUx�;�h��tl�+z��|?�9T9���o������G2��QM�)�𰧳=J�	�A:}U�a�;�M��1|�K���Ӛk����! ��ng
ڇ���V�η���*t����}�R'xG�\ ,��Ϧc�H�^ ]f<�\+�`c�ԡ揢ʵ���]|0�+��k�����L���T�����z�q@�9f}�Ai����.s��(P�t���GЂ���
�)B�<Z.���L#���
�� ��Gm�)}@����g���C�B�� /��7v�oN&��#`�±3���x�5� dԤ���m��j���/R&��_<~p-E91��ehe}�F,��zR`O}Kۯ{��|�f�.�fzԞ4�o(��ʲ�����Rf��m�B��X�g�ղ���"�n5��|��Gd>�*����x�����Y��wk0�.Ő<.g��G���9�5DL.h|i�E'w%J���8�0�P��̶*��;F�����`�T��e�Nխ9���!uR����p{v�qʃ����F?(.:�b:�9�����Ox\�Sm�N��5��DR��^�{+E�<�)�ngx�H�����q��Cւ"b2�`�~m@v����` 'KK��ڧ�%�g'5r���Wlj+//|�����]�+a\i�/q���[QU���� ����.��8��y-���W''��~�^��w�<S�y�PGƕ[�/UE���O٫������z-���k���t�9��6��A|�I��-}���ؼ�� �x'+�X/������Wy���3���ٿ�	�KN���L��5���ݧ�cۈ����sf�%���#�W�f����*����jY��ޟ��6ĳ�ҥ�L��wk�B[Xs(t�u}ljI0�D{v@1�},&�.ށ��ؘ����b)&�A/XEYy�t��E��J�㧆f4�,K&�X3R)p�0ql�V6��nQxx6�l�{Q�"�7b���b	�`P���:�i�E��5�,|���Q��S��`��N&�g�aW�Л�(úXR8���s˸�e�*�z�X�p:ef������97�b[��fF�>����nQ�#�F�0z����G�B��ג���{�����@�تn��?>�τ�3 ���t
O��ܕh|�:[���	�a�ү�A#�����b>�� ���h��o�H�6Д5��i�D�C����篬S��>���%�
�s�����@b���������a�ٖ'P� ��$i$	�'k��⼖O�|a��/4�M��6��)��s/.�Xb�Lb�^I��r���A( �����hZ��w���;+7����Eu����V�4)y,Ϸ���?ȉ
6n���EN�Y�#$h�#�S�j�hB|��l�@s�ۻ��%ؽ-y�:���̩���(iikq'h@-Jt��тd�婫�ьAI%ef�LdL�����s�K��g����!o��3� �H��Z�>NG��K�r�}����u$�� ���K�"���x�'�zq�����das��uv�����, lL�ʫ��6I���9���ʝ�M��q����K?@�o����-�G��ts[L��I�ʥ�tFȧ�^1�"�5��Dfj4�.袸�dp_N}��I�ۣ�������sOI@6@15?�[R����'3��q�� �L~���*XU|�)�y�ש+ĥ�.s_��:�h��S�L4UՅ�=�ڵ{w�9�}���	ME��j A��c�ς��r4oSG-�ǧll�j+��r���(El`м	ŰWDN��_�~6
e�棸�B�Α*�S� ��`q���T$O�#	���d�&�J��kn�Gǽ���Ʀ�����z��\�hS=
���t3��;: W� ,�=�#خ��:H�������dţ/��r�{M��x+N@�XVS�{\D�	V��=�����W �U"/��i����P��0��5�$@tk�~���]�S��L|�W����C��~H����$�$���tzP�b�Y_��8��s0��x)|2T��/"�?���Z)[�"T/;�7T�[R��� ���ڊ�����I�0�{B"�%
� ���/�$-
+P�i��I�U!�V��[�v_�n�����E�4b���0^>�F���Y4M�K/kmՈ&}�x�F��fj�l �4��0�PT�]�3�e�O0�n��Z��^�k������#b�_��,��Sk��k���񙲳ˮ=w��HmR��h?�ܿ��j��9��,��X�&�kM��5�Uđ?466挴��]�ϔ�4ǐ�t��ݩsK$��W%PC-A����?�t�ډ(0�M �t�Xt@��ࢲ�e��w�Lr��ӫ
w�� 5�}�x���%�y�,)Z��q_=`jx�M<|����h#�2	�Gd� h�ªfu���KyV$�k"uS�mό���~���!���ٸ)�t�$�����]�R{�\(�9�g7XӘT���0E��%��w#��"u~�]�NԘ��/�!5y�+=��Y�B��=��>����p�wV.M<��q�Ƈ๹6��?��j�^G�k/����<�!����g|]X�}(����X�fX�qZn;����h�_��	JTp:������S��
�����a-ԇ�[�$�ǳ��ڂ�@ޣY�=�G^pT���,���32�onn�NC�pä��1����[�(�@\փ�ȼ�A~r��	�`l��!�M�b�L�C�̢�_%|�A�;��c!��oLTO܃Q��%��s؈�Vv����PKHH�c��V�);ҥ����f��o�m���$�m�}�&��#i�{ >P��c֓��	�A.\7���5�My���ߢ�E�fɣ݈Vbx�S Z3��T��܃�0V6�5̄��n�{���D��`�|g���*���Vui��e]^��`����.v�.�� 8����~ma��u�gsxC�x�����?�[���D�0�q��K#m7���o��MU% ��%��c;� :�*�7㓹�!�M��S�KhB��r-��G���m�Q���Z(	|A���B�_�x�Ҟ=g�u=�w�~�q[p����e�A�I�d��(���]�f�3�#዗��y5b���|+6���	�`:��	����7�.ҎgD*� q�UZ�i���@6^��/y�Y#�Wrh���p
��.$�D�Yӽ�e����&����jʿ��>�@��T:]p�p_w-�k/��8�T ����7v��*op�ie���d#C�*j+J��\���̬qbg��{C��a�z��Y+ۆ�����W���_:����&I�.P��٠j�I#mi �5������u�W0(�즁������ S]F�u���aށ�P�7���M�2�fp��|v+i4T���_n7��,�%@1��4��~tRKe�U�8BX[��]�z�����`��W��:Tql�Yƽ�(vg4����/�=�,Z-��}�<�7?HDμ�ęn�]	{%����NT.�:>��n���
 �5W�Q�
X��1x��"m�tR�ޟNݗ^J��F��:%V�֬L���]d��Ɨph�-e�"�����BS�"�Є��e�ӌge9rd�R�ްY����c�@�񰥴@��(��x�/�9�S��uK�@� �V�����0����r�䨷�,��b��9��V�KGj�&M�; k��ޡ�܄5��4�L`y.�g������5�#�
��i�7���"���*M��̗�5�6g��UV����`��`��4���N:@�A��꥗
����H,��(�B�ep�.x��>����Q���< ���'�׊N��YM�B|. �k[*$-�^���!�ה_�T[w]���s	��J�ε�7�.lx� *`�	�o�͖y�2�r�(
n��߯�o���W fd�//���Z�>~ l�>���䡴o9#�{�JHƕK�b	`�b?=o�>����������ט�6�v�_�:$�.;��o<(�7�)�R[2GP�!�ve׮]��`v��Y��x:��?�fo�i��h�4�>;o�W����9�H� y�2)�ݣ�] ګ��]'qZ�A����g��7���nm�@��H{�.���ێ;]<$��
^��y
Ի���0=�ӧN�`w"6?����~���7a��Z�!�k��Am�knL`u6@��şf9�J�,�7S�P��L+3�N��  J��E��]�i�y��#����:�ېbd�eT�6�$L���W@�d~]���1�u�M$,փ���WL��R�>��� ��v
z3��ZT����� QkVT�6T$O���n��˂����N�(#"wVL�{S1(�y���P%�G�ȝz���=0m����rg&��_�TO�ih�ȟQ��@��:W�e �$O?l!��A�*��'��c��+&��n�=sb�.ŵ���:ŝ;�ԁ�
B/�M���-�͸���DV�\�>O�,s�Z��,,ۭ�.��V�������ǆ`5�~�^����?�
Em�w�}����Fl����V�twd00�#�-��	-o�2(��IfN=f���H���Wk���C��\U~æY� r�:�j2�Ж���QlBb�Í$����L�0��7��Of������f�����f]�%�z���Zɕ��F>z�����]��P�1ŬO�a�N^��S�4)��u���K#_Y4K�)u���8$�{�~	�Çm {�a�EDD�yx5/dc�j��V�1�?� �J�o���oM�;KD���2�t�? ��H��y��/`sh������b���U�c+hk��)t{&�NT��ei��5��%`�D�oq�Q>��	}b �L�%A�BEr+�s��sQ`B��oa��p/R���KirH!&�����CP���F�d}PC��,��[+�7��J����&���.AA���8�K,��]��,����A����cɂp���x�V�G��C�%��a���c3�-&�Q;�w|�<�s±�pl|�6�O��$b��>��d�U�����^�/�zN���������+��e��Xn�\�M��S񬷠�M���p/�h�]���|����Ӛ��91�?��ı��7��O&O����M��
�1��aU���y���s�c������nb��b�t��w��HUo�歼w;��I]���/;��eܾ]oZ���s�w�p�>�C���O�^�����o޴�CeO���n�d_�H�8�b�:?���V��-X��S�7@�%�>�M۞�ֱ�e.�m"�ᮈ/'3}F:M.�U`���R�gs�@�ۇV\�o}}�O��]-�4Oܳ;F��[�Ө�-Ļ7�iI�Z-!b�T�N���L��Ů����M5;Sz�t�C��e�">kF������?���P�����^0������s˳���1��ؽ��� A|��g���ބ�>(�z�d�V����t?�i�E0,�^�:��SQ�
�^A���Ù^���6��-=-�cm[�� �W=R��G.5QR%��ߛ <=2����k��s��m�j�M�}ὒشѿ¹vxx8�/���^ۺ�0xsySv9e1�5c�֓]���0oAb.S=<lH��ɢ�-��!������?@E���;/_�\{y�u�(��9��/Z&��T�t�=s�E�i3�q^�zzz���C �nO�.J0D~z;2��C�s4���[9�Gj�?�QV�k��"�Ж=jh�����w��WX��k�k�XBػ��6�K�XX�#��r鮲@Fҝ;w��lR?Dus�������NP���%w����VP@����JS���/D�ʱZM��I�#�t��8fM�%���j��0��1�+SQ�:�q麼���]����Ճm�ɔ�y�yU�"�L����'gm{}`=����:��< %!�s���2���9���51;�E�q�g�啾}��n�[���b���p�l�svt�6�J"��}*7���B�>D��Snl!��k�W����;�ֱ��7)��cK�G�����7�ƒ�H��*�!�~?@T7�ڦ\�򩄬��q��wY��6��yDj��M�{�tc؊���=$��� ����py�l�0>�%�ܜ�ajbR�Q�O��Du�������`���M*�"Xe-X�Ӽ���O}�����!��\m�xE��[�wL���gߒGFF�
̉G����$�J�MNN>�:[�Ј�߲^���c��?�-'d+���ӯV%7.���Lp_?y��R��q��Zi��g�
A��K�u��l>g��;���&�
!�\.oR/0Nj�1{��>	1����"!z8�&�.���mdT���D���L+�L�y.�;`P�]�m-荣�?~��v@*K�#L�v�)�w���I��7Щ���+B�g���Ͽ����YQ~�F��9�!��TW9��{����Ǉ���zk���\.�eO;�yYA��>#n�)3��v��V��{IO�5��JNuɱ��ȴ�e�+.+w�[�Vg������.f2��\���i����)�A������@�q|��u5������q��J�٥�	�s'tM��^��]�X#���7?���������I?Z�E��d���D�,��9[�O��A�%���F�Qä��ߩ���!��#��I��?ݹG~=`X��F�Q��4�����==�6!�k]��x7S`��u�VE+N^�VYuu��!��z�0-z�O��h�l��$�A���n�銻;�U�V���^��l0��u��]GZ��j�x��񔁡��C����'�7�o�8 @\ݓ> d�8��9ƉUF:��#�������7�5�A��U�&��[�Bg+�d��΃=�6$��@v7i{MQ�-8@�[G58b�_o��ؠu2vi��6�2W�X�Z�V���ӷg���L�!�˟n>N��j��O��>���h��J1G-��?u��ڮv�̔���q���;RK�d%�ٱ�x��lo����Z'5�F�`���w�h"�����^�¿�����3������mf}���3�q`�r1�����.('��D���FF!dϗ8��󙌜��u)V�B�~ġ�T�Z����q�1_pyjM#b���,���>D�9{��m]Y9�G��>fv����T��} s�i��{��AX-�hi-���������T0�%]�v���=�޵���&���WC���D8L���Ǐ���m!%�_se�����XTi��I��o���%EW�<�u�~�/�s�C���˿����U�X�����t�[� �nlkk��$*𤗖��â�;"K2u�m�s������V�� \�w0�&���������E�:Ւ�W�`
)jkL�ȣ��s�啊ʝ��?\����<DiUp�MÏ'j���]��'m�>}SM=���WR}�z~9}��ɍw+���i�E����c���W8s0�({�^� ��2M��A��
=z2�F�+�ܳo���Hɖ'���+y��XPD����@YY9��Nk��V�y]�@�1�+,�&ɔ/�N�?4I$4�5r��tχ���#C��d@�c��I�o�+��tA6�E�͇�� ֝* �v��z��w"�j��oj@�� �ͺ��Z 3�8�Z?*)������6���K��$��8Ć�>�����꟰����M�j�~>��9�<����Kpp���=w���a�N� �'����v?j7
W{<ٖ{�ں���q���Xn]ط�NI='�d�G��DqP��C��B2����!C!���2g,��%d��92��Z��y�������[���k�u��Z{�+A@�xR%��?�]�`u�ǘ
�7X$�d����
���O'�=�z��!����L:�؟�� gBJ'��qiw���h���q��0��}*ϐ�\�T��>�����P�ē�Z��Wl��w=�Y���G����������mov��D7:^k�p�>��&����۷������ g'r'w���eX��R����N��:	QS�l:g��W)C����bi�xV�;�E+��i�*�B���9�0�
�x׏���6��r<��A7
)�����d}���.��j0��������U2��z���7"��^pb2N�b[�����W��)3�p���V�W&�`�_@��	��S�����1�+���[��~�#��~��=,}���ӀN��4�Z�w��Bl������'�g�&���x��^�v6���#<ˊ�h����'��d��,TW�5�f�a�w�a���_ �5�lZ1}|����U��>`�Mr��)���! ����O�G�<�I�b����9F�%?^^�����67HE�����@��|V�f���M�z�� ��s�A�u�]?�gqq~]��`����}�n�$?������1��Q���[�n�h�+S\�Ad����f�hN�,|���	8��I�A���,9yd9$��">��/NVrF��9��,m��������M��"[~TLH���~b��k�#��J2�
(=.� �#k0���gr������f�<���H���F�ل0^��u�ͦ�j�,77W�d�/�$S�@:D�&��{EĆ�%��z�/���D������-!YVa�A���m`�Ǝ��n䔿��孉��ˀ{�U�KiԈſ�C�U�^�WX;���##�k��e�HfK�wm�/+�<9�'��I�&LD����֮g��c���Iɐ��ЀY��]���#i)�+�Y��,k�k{p![~Y�MI�"�-�0՟����O쑑)��kׇ1͕/V���%�L�x�p��8��o�."�z�࿻ �k�S��jp+��f�5��L�ԗ'�C�>�j���j����)h70<�[�Ա|ZQs��AR�{�to�WS)i���"E2&&&U�OL3��/�v~�3�"d�Q{%�՜��Z4GRu����ł�h�Jp*�3�#fN��m����
�	WI>T�ܝ����G��M^�65������Щ/ �a�k�s[����_�}3�Z,���b���˳
����5B����0A����}��C�i��]h�p�g�㲣]VD�vr��T�/9M�Y�'�J��zD��4�vPݿ�N���=��g��t�(���yyx ����/vPz����+����Ρ��l�,m�$�9w���?��*�Gs�Uh��HAof�U����?#;w��\[�r�ק���ι�M�"ۇ�&ơ�(����R�f����:m�r��־\Y���Z����&����MӦ��O�j�C�i)��z���f�A��}����4jPT�)��.0Okt �m���ѯ�|p/��!�|���
ܜ�WV-o�V%�j�YZckCC�=��I�_���|�m����&�r�=�C��p�Pb�"��vs�̝O,��~����S'a	?�A@X�죎E���/�=�?��T`�F���ԝH�3�#���y�?��1:�LW���}�	+��P@m�}�;9��=6��tkO����d�S�:�%A�ϫ��U����g)�pj���$�W�:��N����:D{!�q�P�=�i\T���3��������P�/�+VsA(W�څ��-<>�A���&������uB��o+G�7���z��=�G�9�0UHϱvEA1��zb�����N��^׽K"%`���>pްc@���٢�z�X�b�DD�\|���}(�C��D�/�m��`�ƪ"��W�����)Ym�F�>�A�r���Wp+����P{#�=��ǎ�kk�����}�/faz��5���v��!ٷĒ	ҕ�HZM/�/=6H)}c�Ƙ�B�$��_�`=�I�2x���e|��@R�y�_pu��ǖ�
UI�ohhK�z7�˅�1��JnZڠ=���E��n���ԕ{�/?9��#�*�	��N����<��2�T��&Ӏf ��x_�����h\����e���\ �q���N�5�b�q9��>1~�j��q�?�P��ZHW�<��o(�8z�Џ����Փx�B𢯯�,*�Ii�鑌�!$��k��W�\Gۀup�y���h\�X�/߾}��Y�JFk�~II�������R�VY=�Co���#�?O�f���Һ������:L^g!��H�%2G��?���ur5�RGW_3Ңq�"�k.Qg`|�x��umD����'/���f1z׾�U��]7���_3��H�p^;�,������\���NQ��m���d4UX����3 �"�lxx|��p����!��p||�K�˦'�4���
��)�R�T<���)��S�l*e`j,G{ڏ�'*�E����*ǯ� 'M�o��d�����ͽ�
�x:e[��X����{��b�~��$���f�{6�S��j�C���?v�B��,&Л������l����>�}q�S�D�\
P��,q×�#U��Hb0�/�!p�'I k#/�ՓA[\tֲ���Đ��D�~��������`);��2f���"�ի��J��{qe�R��Q���u`���lU�z��d�9�7�cY�(D���}��ڹZ4�pq�?�m�WJj�o��S+T|�u���vy�X�A����~���@�Q�|e***Y�����%�R��c�	o��T�~�z��C��,���"5A_�.!��Si����x�n�fi��X/��8+�����X���qn��R�Gaވ/zKhr�x�C5��q�uZ,��뙵lr���/;�܊�E
��,�߆q^mU.
YYUN�X&V(,��G)��n����+�J�e�r~�/�`�IQPbQ����~� Y�R�IF��	ׅ�Xb~�}�C�jw�n�6�.A��S�����Bʔ���@�_���ů�2z7Y���8�-sQz�A�a7��*������"u:�Id���O
�v��j��E�Y��^��� 9�?u����#�-��ªA1ovf��a�F�Vx�g�n��S�x⦖����Пl,���i>ߴB�MV'.�!)w�6�d+�����IX�����ԑzSJ# ���M�5�SX�||'�5l��NT+��db}�~�eF���˿���"�y��2�.��m��ͯ�ƀ�+�j�K��¦n�M=����b�f�����5Pߔ�
U���
���NcǾIi��Tj���Wǻ�3���ч���������W7B�� �R�%g E�Kv-��'y4CVc ٢/��r"=fi��:010�{�u��9j�oo.��cSʂ4�n\v_�6<<\�:掶�}�a bPhjj*�,4���R���ܛ=�<�1]��=z�g@���S��I�
��{�8�{q�5א�5-� ��}�S\��o�o�/	?--Ř�M�%%�Q���H�����0�B��"��ώ�������;����&WYBmw��P"��v��Wp@���8~	N��g:��D�ʗ�q�OW�Kv�.�7�%�l�x<�Zw�5��qU������v��n=F	
r�Վi���9I�'-���?��3JP��<�w���J��}e��gŨS̳��C�"���^'k3|L�M:�������h	[~��Ǧm�ݵ�F�%���� ݄`��������9���~�Z�oFne��<&&&�����zE+����r(M���i}��Z�g��CƓ�Ȉ`�����\��}`�M'?����j~��)&D�t��ӆ�_��D�q'�R������>؉���~��)���ȿ��~��R�O+Rw粣���=���?���B��9�<CZY��3f�� ��^����R2�[P"pj��ŒL$�}�A[��l#����b�����O�.�g�n����|�V�B�p��"��5R��r˔��&]ՠ"�N�/��}�'�"R��'�'�-����G��Y4�BD� Yw���)�'o�xE�]�O��v���]>��B�/V0�M\�'�2���������v4�v��:��mI�B$m9��R#�`�D���������Ќs+�#��?��
�W���R�ΐ�#��$�4�u�Lƣ�{���
x��/0��w�O�	{����-֣\,��>��˥��+�/yȼ>�i�����'k	�=�D8$�� �<��?2b
/� m5�jO<93���ۥ8�(U�/C"���C �%g�OC<�~�]�9��6��僫���mbA�|��l\\��ec9r��������d�1.C�ڪT?�G�#q����j����EX6�T���w�E�z�H��gj� )�|a�64�_�Ʊc�[����{^��O�I�e�Au3���9��eђ6���]���i��C"��	��ov���������ĉ����0@�/���9��X��*	"�P@��.���،��mJ>~�h@��V� S�~��-�]�#����+d»EП���F�ʛ�*�`r^u���2�췰8EۥZ3>�\� ȥ���p0ƿ�$���/^�5XBer �A��>,M{�V��]s(Y��`{/O��l����p���D�}����ܘ?�p�mP�٭T�� ��X
d��Z���P�2����P>�9Y{�!��y�M"W��Ī��n=�Erk����[3����}8�֨YW1hFqI%W��:zd	�O/'��}wV�Xl�D�	v�ky��Ƥ-�''�h��[T!���N>��8��T��@,�`-Ӈ�d����*!Z4��8q��vI�a���"�r��i������+�h v??�������'n���k�����W�g1B��U�D]�
���5_�}4
�&�(j�	.��oF�% ���7Q�D*�`��\s�N؁� 4�o�S:�y�?$ݬyn�T��Ȫrѯ��oԀ-Z�P�Cv��,�Q#�Շ��A2����ߓ��/;���`(��92�Ǔ���:����_2���r!M�W�ȟ�'�Jv������oEz�����<�ڸ�xb���---���:�A���O��K�Y�r7I�Ȅ
��η�9 ��Y��(D���$x� �u��^�C6��BpcS�(o�������i�ErN���j���/�}�ÎXˬ����NQ�%}�y�7i@��w_lC�!������m�ԝ��L�C�?7Q�$�M��w? �1��U���i�Z�O�flb�!	�����W��(,�\x���rk둶b�rϿ
�w._V���%�9�ޤ JMƳ ��)`<�#�����4"���M�Ż��?M�D�qƹ㦓oI>YĔ������6T�g�A��rL��0QG�1����@�~ʕ�@��t�d�`r�g.�&՚%Rճp�c⣷�w[��N�8P
�1#N�Kb43�dDD�qdR�N�J��o"T/�ju+|�G_�h�3K�	�Meo���̇�t����ӿ�M�����2%W\�W�%�l�o!{`
���Vm*��F�E��,��a{v�頵Dc�}����vL���x�OU��8	Nk
����W�ʝ�fiƓ�����2��E)�`L�X:^2|�lD*��a�v��w�~�B������L�&	��@���^�Uu��X�x�6�'�U�e�jPN-�cנѾHy�0��P�K�yNw�>�ڄw��꜁��nZ���PrX���4��	Ђ'j3�~������a��m� H�S���a3A%B
u�\]+������+�ݻ�S%���yZc�#�7͵�X����j&�����?u@Y[1|˧�<��jV7��d5����yŵ�:�p����VY=���Ո�wV����-�,�;B�|������ghu�I�kW���}� h��u�RGA�D0v���!))Wk�J��ܠ��U�A�i�k�ڋO>��?�K���kI'�=�-.���v�C���j���x��l�9�!����G=X%S��k���Q�����G�*�2�WT�D��>��n�U�����4�?���T��h��8I����Z/v
�Et��؞[�O�B]���/..އ-'���ߥN�E��[H����Vۏ\����t��> ���u$ٴs�h�Cd�y��'�`�T=�I4�Z��p-G�ip+A0�G�^�oZJ�I4H���%���X��,��;��K$p���Y�>0�̭]q��-oo�A`�Φ�x,�,��:y�ONS�Hlц/ҽu��������e��=�Ɋ�a�8���5�����c��:��79:	-�-��%���b[�|�]b���v7I�`��{�/�q�'�R)���������&�E�Y���:e�kk^0䛘a����	N��g�{j��1���[���~|����xx��뉈k�b���r������0~��_�_&��"�'7�;���-h�o������:��:�n9�S�[���_��C���}���:n�^ K�� ~�ۆB �C���VTD��O�TӮ"�X�\=R&��.6�:��&�i�+�
)�2~Ư*E/}Z����Z�&��u�Ux�5@yţ���o�_&pG�&�Pxx��@���@]��`k����sk	��|�j�Z
���ǇXɼfD����������]0/���$ԲӺ�3s����kؠn���Ǽ~�3�N�e{�����m��a;�t\�9_֚Yb-��hp.�S�X��4'V���y< ���;�y\��f�� z^��@����+�|�~� lF�������I��PXX�8I~ r�$%��,^�Yn�V�0Dsb�\\5�V���^�P��'s��Mh��-��W�!	l���^�,����-�۫������϶���g�4h����g	�`+��Z�@����D��;�v��yS�|xs���lњ�:�` ���6��SYYY����Q�-���.Q$�3.��x�g�b9���s`��F�oI���N�<���	�"��l�����t�����"�,�9�V*U�<��)�#^�'��2 eN��(�'O4�9���w?��]7�o�i���;E�G
���wp�2 ��g`�3�p�|8��R=f�1p9����2y���ר酸��0�<��B��|׆@�Ҁ�oI��O^?8��ԁ�6���_��2���Z�y�UJ��}׋���'6��ss�As��. )z�'�a7��l����r���DTl���x�!_J@k��c{�p�g+����x����
^<��h&���M�!/�>�`��������������ϊq��8����KG){?���0��� B�����L9l�6�����ː���s��ţ������f�F��}���t��Ej��Z�!��.�8�	�Yꚛ��FBq������B�Y�}>d������MB$�עiI$	�V&mݚS�t��N	��-�g��)���>�U�0�3�\�FS;��܈�����G��F1��ƊP�b����Z�ڍ�w,J�n�����V���d.Xf�Yy���䤧̀y��N|��'exI��6� ���g�>�w���P#�5#��0
g��d^;�n��G\��������
b�wq%/H�I���h�%�?�n��yL�L��_H�m��p ��m��!�as��N�p��|����y!�y���eMMMo�ƌ6X�i�D��
߼pߟ4XHkO�#`+w�3���`ӆ3����u�T�y�U75����m��;&��%[�J`���2��,5�-#�G��`�o�^Iޜ�����8�eJ�����R��D���������q�J�MUeew`2y66~D5膀�+Я�̃g^���v��>ò�J��!N�\�ܢĩ�̭��&���HQ���ލ������$�#:�\�U=c@��lւC�<��������'͡?w�ۣ�|w�QW����¦c��h����Z'�C�Q�O2On���0l��$�LS��5���/��թ�U~Z���C2%+� .�h}GXASb��n��H�K�&V�^>~�GGǬxO��$��c>;���� �czH5H޼�6ޛD�K��">
���%���Bo�H25��/+��^A^�>y�k�y��mvv��@k7�=d�
�&�r�ib~��R�F �O�D��]�ғ� ��e�@s�P&��Ģ���~iJ8^�������mƛv�W�^��w�2�D��UI�OL��Y퇻�o���ln2��0��������� !�$����+ �8���[U�nW�MR�Q�VV��w�
��"T���p��BZhH`Y{=���y�aGN:x3������&ĐΜ����*N^�%�(��rf(�3�(fIh��7YR�o!�0M��,�u,�i=�/��E�l�����?).�d��@;���'�i��%�������Z�k��1�w�h�B���mҞ��\%��l�?��M qȌ vpQoR���|de�^ԋ�9sbU�Γ(��E9OӺٙZF~�U��ׁ���߿�F���/h�����4���
�gX�W���$1�uݭW�澞��qxƼD*�ҥ��:��u�2��:��;��W��7���]�(�LD�}�c�����+�%������͜��Vŵ�1L_�=�J�h�ecFj�~,��~t�ݹ��ˎ�����ʃg�Z�k>|zy��q!��{x�\�Ĭ����Ȇ�j�@�y�������vhǽ�U�V��г�eG)����>魪�;���`�ׁ��R.��L�`�X��,�#�[�>.����B�QR��V]]M���b	��{ʪ��0����HPw���n�jx���@^O2�;x���{�k7?��#��g��%������Q�>x�h]l|�F�8Ԕ�^����N�k�qgf�VHp�]�'�<)�̬>Қ;�K�ACC�C�扩Gj=6#8	LO��v"~8{sx%�Q���{PU���;��)�Ma?��'��N��FX	H���.C�4�	Ss���;�4}����+(Y���Z7+�A�����/0������ZY��;�4o!��gw-�v�]
z����9�tH�;"Ov�,a�ٲ���������6�~�lo\���'���o��j$�����<����\��)�� ��f����.>�>v�M��)81Ծ��C[U��OW�C�Y#Ng7T�ՙ��F��3�l[���>����#^�T=��74T�����`p�����p[��oʡ���WGX88L�ad�
>jYV�l6jǎG(��w�u��F��>��  �xȑ�P�>Ԕ�d�ϗ����E�|��'��¾$S;/SF?㯡V����z�����ޘY������?v�&��'�^����{%�����W���]Ğ���#��V(�/�j,/��N�^�nY�\�u����b��^�nm+�k=^F�n[��|g����of������r��r�/+��E���FB�Z������MC���ƴ��*"�{ӆ�����[%m�5��sy�S=7e��+N��|;��H,�~�������xl2�lp�5.�sv5��M�O�z#L���59�&��(�<�~�ݑ������q�_�#{j�X��(�l�*����̮�e����-��ؕ7ݙ�pV�_����kXM�GݻwO1�B��m����%)�\�lV|8_�w���_䕏I���s��[����T ���o����e뺊���HN0��B�,Qw��_��a������1s���7]�z�񊲕#�.��?��C�>��D�M�R�-vN���a,Wsݦ8Fx���-�݆j.-�R�"C��U9������~�]2�E��ǈ�LL�H�ѧ��}���i��2�4�#���(��WQQq�.|`���Q���q�ĬW�2i:�Mg��j��l[K���b1��1�����ѼJ7�u]Mߕ��\�Tt��-|�C~�.�����gg��M)���������
��[%l�O�B���a�P֔�CN�L��c��.x֡V{e4��^���FMԚ�-�C��3�g`5�\��sqɂ!�n.���`@ۗ���K�/��N��l�x:�bƏ1=K�$9l��/ W�r���Tw�wH.e���ϡ�T�m֠������Ne�=�xt����:|��ޣ����ɳ,;�:ɪ���M�����EF}�1��Â��)�D��v;��$�X�������LVuZ\ͨA��2䨨i�C�/+�p/Ӑi����V�Ǎ�ljMsw��F|���+��-��s�%'bh�`@r�A��T˒�f1]����Nw͝���ˇQ��'�h�Vv�8�:r�o�!����H�6���.����>I�8�������*]��8���w94�*�.E]<FFb��( � gr�Hc�s��f:��"������w8�$TKC�?��,��f��1�i���܂p� !�;�X���;V�ׁ1���sn�b�:~���q��L�f	s�����62��_N�,�KV�?��֡��B��<i�/}WHTRI�hg�=�W���~�~�~_�@��S0R`YJQ��D�gyO{�E9����h��p�������"�rQ=�dG���_�0at�_�}z�����Mn�.��@uR)RF@����J®��S��db7�\kў[g%|"��ua~~��N���b7c�I�tU�G����&�E�����Z���I| @"�2���u0�S_Y�E�]���ٴ�����a���(���|A�r5�6���r���F}�b1��w����E{ى0e�>
���}I�O�v�vj�m����m�1h	�����Բ��?��fі���p�g�`�nff��/�����¢;�a�6�ք�V��7ׂ�}>i�?���ĝ�M�p�؞�A��;L�'�e�v�)#H�>Z���7�iu�veb 0� ElS)
'_�M�X8B��﵅jU�z\��3�&�� e�(��PN����
�+��Я�S�f^�Z���?��mdʺ
̒�b��������O�T:��"{��jj���#w�ү3{y���V9�5����Pϰ.�V�� ǇZ�~�j�G���5�، 0[��;���u�k�����j���M�X9�P�	 j��x=<'���o&�`�<�����R�4�M)��CGD�(�͆�*��
�:�4>��c�GǏ����>��|ט�˻��0�G������>�rգ��a����#N�z�~��mD�H��֣H��D�At��Y�X��V-��`���C�փW�U�� �������y��p�>�6l+���7$��{�&@J^���ħ)��9i�P++��k��BZ	>��j�O�= ^}�i㥈3U�A���e yA��q6o�r	�gN�
�S(����i�:���)�����*�ÊȘ�h�^&�1�s�zdC�"���(i����2�q�c�����q5� �؜I|�����e�����e�")�8��V�ЯN_q�2.�h=��^墍��g�G��)��c�eb�ూϦ�߀�<�kj�T��S�%?7�8<r�q5g���Ϧ_�W��5��hr�"�c���$��W�yt' L1�=�>�����ؠ\D��������o�6E\�K���[4�� [��Us�����b���c�D��i�A�	e�S>EX< &0˘�ĘyP8~mpE�����ٯۛ%r?A��>�u����m��w큔ѻ�Ad�5A�F_0/��x�Ӿ6�
�L)�@����v��
"ux9�vƞ������K.�����.]_���jY���JLvJ��*��|c*-�D?�/&�n��q�E	�8|�:�u���4�pK7�.U�"sQ�PZ�P�7�"�Y��?�oW���]Yb8��+O�rl[+`B}Ssq*E|ضH��ӝ&q;;0�P���'Z�2$�'!aB>��2T�5��&�����U%�;M���߭W6~,��{�v��|�+[�\�Ӭ�,ZQ�r��d��˷�(4�[����~���@͆���Y�~��x�/0�����ö���B �q���JH�A(��3�X�G��[?�|��,e���CO���t��a�`U��o��D/�����
X:�ġuBZ���gr���ޅVK��É�]�!8� v����죪!������.j'�a��6�J�4���!���늚h�F�����V������|�k*)9����i�~d*��z\��tV���&
�gi/M�׋m%��u&�ieW�� 	�k\�M�}X��*+G�CC��fE��\J���i�tqll��>��l��X&��#�M����N����n�]`��&.�i��:�F6��=�aq�`(� ����<n�`�RB���Ԝ�#�M7ɷ���s�|ku�o��_��� * v��ady��ի�K�奁���P\o,C$��8w���M7�	�e4��h���T�,��{/?�x=De���x��={'��
���*_/�_D�������^�$;�5᚛�U?���q�k���|� �7S0_i�M��r|m�'��n��ی8|��v!�lv�6�'��+%(iu&&2����;����+��#|���:�72�1�惼��!��6~��C��-[bˏ+��_U�	 ��� �餴N�49�pLr)�U���G������>j�/����ߨ�`������~�q|���#G�(^�?
~t�� ���ھM`p��0a�L�_:��U�i��i���7�F�L���#���!����և�ԨMa'�݂5Ƹ+�r�U�/�ؘ<�� �f5�,Z{Yp��P�P�|��&�
�9�ǩ^<Ŕp����G�JSJ�&��9�2Lp�p�M��Ʃʪ*C�R/�+���h�H�6nʰ^��Ǯ9�W���{I�(��i���t�Ѷ�hz0���P��W�[���<;`�𙷂|]�,	�~����.�5g�2�5��P���h_���n1>�|��� `�W�����J�qW�	�#�3??�n6�)��
�Crc�b<l�CvK}�~��Q;�0�H�t,xʏ���ه�.�M)�(��g����n���$�֘��/S���X@(577��HU3�#����	��l߄�5 �9�O�[��|�R���' ��������f�ܺ7a�� �
 ���Sǔ������+�n���FpƏ�V}��KA��荫r�1u�y���m�*ii�	�R�����a!�3l��2	D0>n|R`������Ν��W�:�ດV�������&�Y~���2<�\ĳ�4�3���� �as����p����9��f<�0q�����VxI��v�Q���?A($�x�'��94M5E���S��Ņ��^r*���ы�:*����Egps����u�@���!Q�ᆻ���eg)P�,uC,��"J���)�w/�߾um�O���G���jcZݟ�^&l�����1Q���*J>�F��T(�r�ۯ���m������=t�	x	S��W�o�`�8_��Eķ��;[Y߂��^�MEӦ��� ʘ���O�1k+�X���=>�hB{Z^t7�����gWs����Ǌ/��#��3C��CY�I�#���Sy�V�M�6�_K%����'y��5�f��۰�)�a!2�2	'ky����[��t���8�]���X���H�n�M�+yY���R����>\QQ���L�+{A/���<A7��/�*��/�^�;qiiqa�hl�.�w|$�2�d�ˣq��p)�JD�!�<����L���5�����/,@>�n��*ڳ���qż���_B�[3>�ؐ�K�˴����tt�����u�#�o�b;�a�`q���M���O�-X6l�i�r�3�~n(#+UWUҊ#��u������X
8�""�Nоb^5Q|:���V�eZ]��M#G�y>�9 ���GE�o��a)m'�c��cX5����-�c!��Nq���Dy�I��t�ޅÃ\	�� 	�}G�g��dAn �s �8�ƺ���L+`L��]�j��PjM%��ĥn.�_I<��Ue�NZ�&&��IX��3�Y:2k�+���Ha��S�'X�h�� 8F]�gS\�p��q���P[h[P�����Y��[��,�8�O�.��]�Q	P�Е: B?�a�-�N)����5
FO���t1����ծ�4 l��? ��)(>�)�"/ʷ�"�m�~�=<*jɏ��/9uV� ����n�*�6?�-�oct��݋mv9��U0���2e�<Ho�X.������!Al���q�F׻D�+D�Z$zp�$�	`�U x�qc
�]��� �mA,(��aGj-���NFԏ]�kY���v�Z<ʬ�/�!L������I���X\y%vL.&ڟ���wnr�͈&���?<`8ܚ;W�Zp�)˾�3��4Fٱ���	��]�b �������w����[���H�<&�3�Vg��Q�oBM�����	�r�����Q=7��<熰#j�1�l.VA�+:��XC��.���,����㊡s해�ʺ��^{ѯ�����j�f�¸cd��s�!�p�����S;v��y>�*��<�������Ç�<_����绐});_�T�B�ی�W�3��ʞ{Z�*<��u?��W������ RC��+je��j�I4��U�|sd�}G-���{�yx�џ���m
2X�M�I��*|\��p�}�">�mJA_EN�%°��zsG����X�(|���	8��ESim�z6�5X�?~ �x��H�	�h��`�Ƣ��F*�~{�='�8+&��׻�I���L��Wӗ�	�Z��8����;�n���D�0����(�$F�m>��ӄT��V�����+�l�.c=�\W���݋*�g`j>�w(�װ���hϚ#�����cT��Df�S�/,D��
�X`�"�*x���tDR��� �V���=:�梇]�F�>���aw�v�2�#b0�-�5mޞt��D�vt���6�ߔG���* G�j̰nӭ���oZ�w�����q�M�����L�q�6 �K2�]����XW��\�A�V��hʕƽ�t_ y�uoc�ꝇK,�09<�*P�d�S�&U`z����i�LH������lp�8�������#I��Ċu�/��
a�BT��O;���8�¹�*{���|���rd ,���	9l�EH�|֞����-�9_��T�<s�XMMĆl8\��l�SoI�6rdP�n��*hᡀ ��v�Lh[K��\��	��1�0�|G���2�]埜 ����\Βd��L%k.:��߀�h��MBB{���C������v��6���Td��$��z�]6��9)�� R�-�J�~\auU.�b[�ǚ�i�Z�rL�g�P$�\��`�awk�qv�o�;���<�_�v��=����D�W}7O��l/�:w�[���y�e0s0�(�Ѥy���H�,�S�N���U�f�Ȯ0+�_�8qcچD	��=�i�A���hχs8��{wI�an����("X��qs;�pO2����4�h
��bBڣ��a?8]�)!�w����NV���R���6R ~�)�P�����L{-�����Dw`����@�d�fn��#+}=��¯����װ���涚��������[��o��4`��:l�E{�)�2u�L��\�@XF����ͨ����v���L%c�
������4�ه���3|��&y%?WU%׹I�L��òC?(�m`��Z�������*El �
4i�}k�u�oba�[�b�8R=O��`��U�!#�[/;�1�-!�Wq�K��!���a&��d:���g�@�R��<�j�i����b���Ķ8�a>�=OeG��]��\�������	�Fhh��f96�٧�P�ſ)��_3Y�r��4�WLU$$$�`VK奫RT�3��(���}�n�%'	9p�]��9�H��7
"+�����إ�ļ�f#ѻ�`��iE�R�G9yAEQ��񌦅�� ���-�)�� ������'�tu�:���YGi���a�ػKLl���4���[X����-���c�G����v�%�!�<;\�rj�
"�3�E{(�b͹Z�]��a2�%>Tb��w��	���7F�-ڹ��v���#�`��lmG��ȡ����^��u��?�9�]��XڇϺ��3Q.*ĵ&�,ż���:~�1]i�AM4@����H������v����2��;$Ꚋ��촷ogo0x �m����a�@��0c46ُ�_�C������B׍d�nC��M�wsIt��ٺj3}�M�a���Y�����{�6�,�Ȋ�gOL�!��1'�a�l-�9W5t�=����5���P�f�O���u˄߫������k�ҳP'��9+X�y�M��)��@��*���l}��{2�� �!𚚄;%��"�"�I�аx�K\k�`�����9]��Y`��xl'�p����>y���(���ጝ����Sڢ@vgMw��S;��{ݾ-.�	�� �\�����D�b�����6�����~�mZ[f{����#�%D�Qi֭���?}�?�Y��P�	G�<m�7K��Ad�ǆx�PW��T0A���h��P^
���/�b����_.}V�C�j�����-�*t�F_�G5���B�<�p�R��zN`�Ġ��ϼ��Q(�G������X�]���{�6䈝^a>��Aw�)�j��SL�;����U?��d3���z� >�.)�
�8��gp-��g0N�:����)u�Y��yFN�|/��9l�dC;���t����=pb��2�D��"`F@%df�����uhi=ў�Ϧ���@2O�=�q�6�K�(���{�������|ɽ��<�Y��j�-ķ+iu����@��i,b�J��#ys�X��gw���H�rɧb������
��v.�k>���Ν9r���e�U�D;��k���g\�/�2Y@֦@�E̤���t��BCV�/7sX����Ut6$����yG���5Ӆ;��Q������qH�v8f+�S�����)N��K��c>���l"?~�o�?���{/Ab�ݬ��bO\+�T��f�b�h���d-N�����}�.������������__�����k�&RF�	�L2`�w�f��}VN����W�~�i�L�q�C�tut<%���@.�L�����m/g���m#Q
�^S+���a��즡E+�i��������OϪ�=)��p�&�#L��W,�<YKJ�=���_��V���'��ژ�Q�~ɇ�������Ϸ2��$�H��8������ `a�V�,�M�r�J�k}�H�W�1�El���+�1K�5V�pa�����Ao��R����p;'�,ړ���g��@�:�{8��9�n�2��z|0�����(��d�DEY�C�-�.¼K������.�a�i�f����3�W[���N�����ܔ�`ç'.c=w����)|E>I��-r�6C�@Jʡ0~�a�6��-�����Q)�Iɽk.ߜ��E�3ρ��a�}�j/(��CF�K��o��r�
��*4��\F��q!cG �q\|���O�p��]��?Ɔ,5L��d'�,�rn�����|k� �fk�� ik�O��b<M��oS|��>�رwS���i
.��u\|�u�mV��(�+pd3�������6��K�j�_�d{&�Yp�&����΃[�olNw�a�<���f?�v{ج�ɔi6���qў�5���U�~/�����f�.v:=g:�'J�;���tԑ ���g,-��f��i4Z\�l���L��]�����Z���oy�K��
L�i9&�Ŗ�Rډi���.�!x��^>Zt{������\FeU��y翌��ۿ���oS�}��� ���V)Z�X�]���ܔ�m:M����fD����r�iΒ,�Gt�4��ǐK����r�s.Rt�m�X�N���;��CQ��zB�1����P������ND{&^t�D]��9�oX��>PgAǰV�1aB�v����������3����x�f���J�DJ�g��9���1]266f��.%�m$�7�E�Q�MåP�� ��ӿ`������	I�%\�6f�h��x)�ZK��H���W�#4yr������Ct�b�C�%��10����$w� Y�%(��ə��9����/d�4���NYW�����Ju�u��1���\?
v��4 cI���Q����{l��3�Y�,J4ў~�x,E)E�hU�x�#���"�[�9f0֠��"�R]��`�[�Uc�fl;Qf�8�qQ�-��I���h2g�_�ԯ�
(�O�����!s�#��0!9@��,�ȜRJ����+o3"`��/C���?B��x��>/�o�O��$�)i����/#Sge8�uW������t�=́�Id��[�&��\w�4\KY
kYVm�a�wa(�4�J$�7��Ƥ�ٷiii#�����.��F��$��2�g�GL� |i��j�d�S ���[�s��S�B�J)��$y�7��ucfU�g~�%�^�̂���
����^;��!�7��,�%i�}X���.ů�����-Xt1[RFG����4�����C���KZ1�F��VH��gff�۰�l��5D�# �+�ITl&��ؑ���^��m�/�CƦa�eo���"�Θ�`�);k�ӧݰJ��ڲHe�}�,�)Q ��ֺ��@��"�Z@D�@4k�����q��c[U��a��#��pw(�����4�|���+]E�(���q<�������	�\/�Xw����ᇶI�Rp��@
��>t��EZ��Hk�o�懐\6:4Yf,�0�O9r(��Nݑ��|�wh�C�j{Fr��6����/u�>��"ND��&#�ã	�C9�f�E;�f�jS��:��� }�������C�Q}H�k?�]���ѓ��B(هh�g�ډى����W0 ��bu��_M����-�nK�D�v�^X�VwB]l2D��YVp2d���	�S�	i��Y>�s9E�4�>,�M� �s@��k�z�&�3�&�%�	����&jsZݗ�+�aX[KH����T����EMb�Ђ�k���BQd�Ï�U)�MEv��Ԕ[�i�eO��J��+�-"�µ�I�e���s{������}=_��y��8��y.��RC��K�ݯ��ܹ~�_d�;m��9�'xg)������Sw�����i3O��>Ӏ��dX<c?�� ���,n}�����F_�1ڱ������1�,j����O������ĭ����Zȟ�� `�Wb��7 @L*�+Zb���4����Ԃ��q]7� <�?~Ïk�{s�MEI�/��1eOB�ƫ���c�\�[w�
񚰮YINM�uq����ڱ��$�ؼp��Ɨ���}��T�SǟN��iM��m���'D�������~�4_\>��USU�4���H�U��(8���%\�X	̚Y�X9��,� F��,5A/��on�l~%�z;�2�j����p����y��\�<)�w����|p��X�g�c����{� Uڸ����/=��M<�"D2���7��Ԁ��H ����: �;�]L��:�g)"�]�U7��B6!�c2LU㪳!�t�8Bw���%A;w�� W�3��O�`�+S�p� �����7	�	m_��.n�$��kݥ�6l���t]H*���L�a��
�x���"��XS�;|E��}���8%l�9[��hFaz��9F1.�Yyq���\UX���a*y�K���IcR펍���|��a�2����cC�ƶKr�f�!��1;�=�TE�b��N�B��yY\�o�j;(4Cq���ٲ
%I��&�����u ^�G�(�:�ښ!��1n
T�$�a�#.�a�SBB�p7n��%��{�j�K����?�6W�����ڲ��!���&J����I��tQ��'S��B�X#?w@�+k�z���BF��e[�M���M�E۞V�ꕵ�苩7��4�����Ma��q�`�����h�M�5"��9*��Fǯ�eeM��i#��
�^�80�0��`��N�����YQ�T����wBǊ��57"`��+*|}�S�(n ��t��Ь���5g2������&\�h�S�ri�"�\<��8��3�ρ��*4K��N���ySq�,��Ω������jV��>�р�
�A�9T�sϘ����� rp�+��0S�Ԗ�66F��E���=@�j1�e����	9��3��;   z�/wi��Ϳ���˃���0䝳���A���n���It ���5����Q4���Xu��E,�5��'�' �ZƏ�����}M�{�B�dP;�+r��w��Į�Z�a����f ���Zդ^��!����ᩓ5�����~�_�CKr��f;u6-~�����Rx�)<6��eq�:��ؽZ���#�]�L�М~�B�o9\K7�cՄ���;�����{���#_��q�O]�X�����-8�IղKLJe2�tara�"i�ם�f$��88�\h2�*�3��l�D�����m�[�\�I��7a_��y��9~=`�x�}�4:UZ@y	�
�\�q���V��KgXS����N�H����+�̨`�з��;0�~�755��wǽ����D�'�5���?�%s��O:G�AΊ}e��y���K~sA���1�Jw�Ahf*N�d3"-g?�r�?#��@p|=���4��(�c��B������,���Z~:s���&��ZgS���ťծ�p��߼ySa�
hH�ѐ&I�׫m�O� |�.�7���
cȯ.��p��[�]���
9@�[:#+��O�m�Cx��M�,��:
(J3h}�@��G�'������"�������)o0��m��� �Ơ"�iގ8��QD�$�C�l"��}h��dxj+c,�Z��&@\�|���1[f���d�y_�����P�K�u���6o��WT�v�{�]�������'�(��:�(2���E�� a��߷b=z��c��B��r�&QZ��름k�~hRrt��Zl/\D[�}�ɶ?Ο�[E+ڿ���I�5�g,U/���V��+R.p������K��|=�|(���%P撟�k!٤�yc���������������O\�Ӻ���b)�2N��t�H��pw+�Z�y��;GW�qp�*qa�W�z'�SrGvC��V[h�� �K�'��tuu��K_A"g�+&��?D~���3���טli3d����b6"zO�t)I��j�?4��6qJ�a��h��}k��V�u�������`P��黬!os��mO�#B\QzzG�"~�F����󙌫��<����C�Z�������H�">
�
^�lw.r/n���� �=��$ڟ�^�_
(,!����Ƽv`'WXF�9�����W��Ĝ��6(���_��u�$_ݵ�4\ס~�-�/1Ʊ�A�{ᑋY��Հ1��S�O��QS�A*��*�_ &8����n�
z	��B�hDhv�Yy�=}��rh�a�O�R��ttå�B��~$3��1qq�u�E8my?⸨���Im^���`�n'�@�촁�+�-6FQ��H}wO�3���t��b=�;t��ߝ ����:�v�v���Ut!v!���&�;cB�b�����5����������W^
�| FQ#A�YF+L�"�_@�h��$��j �<�W�{zyO��}}�7����JqW��8@�+�/�.��a��c���w;*2T[ʹ���u�=e��s���G����$v�`���s���A�ޮ
�sF��r"�*\TlR�<FY��|%�D`�����z�	xЛ0��d��X� �G�C�>e��}�� ��_��[xT�j�h)S� � 
Yl�/��rJSS����]�6]{Hdֲ=�5 *Q�!�p�q�6�m��o'2y���q���|Uە��꾝�ksN�0��n����صGNn��k�+�9�P˟`��3�V�i.؅�l��m�+g2p�k�O�BD�)��xp�8j]bNYO�������khh؝!�R,�BVQU5w;i����G�4�`�W�]�[�\��vyD�P�.�ͽ1�8֥��j��_&����|Ԁ�M�%p���{����Ԓٌ�l��`��/�)EҷM?g/������L~8�)I�Pm0)����b�3�ϧ�=��K��2CCh�)f�a��')2�MARQB.��w�ͬ��`]g���6��-3�Op�y�U9���Ou�}��L�5�[j�-���!E����"%��p�#�����Xvj"�;?��[�ȼ�+GpA����}��>+��5F�r�r����Td��e�;�ՠ�
��F��e{~�6һ�DPRw�jɄ���ԅ,�O�!h��(�5�n�C*.I8yg*8w��m��=0���T� �!j�@G��*��	V�C��ܪ���t���۔�N��H�
nܸ#�SFz�Y\�z��	ͤ�곴�%r�! �[╕�j׷����.*�z޾ p�9��ggM���<��n��ҢX�	j��.?����}�1��=���HNN��.�C[�x{�%[,�E�BW�N��:<��4�z��`aI��b�%�dP����:nf2{�Z�a婿[h��H[�� Z?�C��{��m
��Ox&��p��&�`�Bʅ �[vY�����Y��Z������=�\�&DL�E�t��.�q5�7��/���A~�ߡ;U@��(o�"@�,�ﴛ3(7��b$^��Xv��0z��|9H�˞�����aa���_�m>���&�0������]z��WɌ0��J�k g5I�M��Hm��[�鍐.�s* �ˈ�_%4�.H�,�K�C��H&��@M��;�	y�=[oҩ���'_�.K5��ג*d2���>��ٱ����L��#͑��D�丠�v�^"m\$H����ԉM�	�-:�@��|I�Kl�=�sir��0|�C��/j��AW�R��΅Ƞ;����8�=��t�D���g���l�Tܿđ\p"S�{�,.?�C����[�E��]M��NstL���o �VS�]R����1W�V��f��7���(�a��ꒋx���}��m�Uo� ?У��ǜ�1:>~��y�l:���<����:B�6VVVr
�a��S,da��e�Ux2���`�B@Ξ�g�?�	u�rh|���:o�vl��@��W�9�6�j(��BW�t���<xo%Ze��@v|Ι)���m�������rkH�Wy]~{���K��Wқ�}k�Z��S�T��t\Ѡ��p#i�J�_��ȹݽ��w��b\)"��M�g�P�^8��S�hK
(\��cɁ{GRw��\z��=���!�c��������n��b��2��8��6%��H�,:5���H[��-��1��U+����@-�8�;�ї��wR�������X�X�~�4
�<��\w��Ţ�`����zcV[i{���*\oӳg�.k/&��0��Z���q�]��=��g��yά�灓zc�o�\'+O<�l�J\��%�ң��<J?�Kd\��n|
�Ӫk� ��</�_�����!B�����wkD�+w��ʑ��Ǉ�X��S�g���}3L�D�ThJ��S�#��,�d���a��+�H��M
U1�:5��+7 ܙ����g����y :���X�p@U�R�L�_�]ۮ�3���6+� :�0+�Ӱ�]�;�3��&a��5Y�9�i��ͭ��������1|�7o޼�+y�E�ݨ\m����wa���;�����~�xZ����G[ɢwi�Ϥr�K�̮#��6*s9�!E���`��9�ӽ�j�T��M���H�"���Աy	�BD�p�e�;̶CD��q� j�z�XZ��>��G��q���}x:.�����Z�e�_�$.��o�Iu��ڝC�:��8����´w� a3�)W�o p[k3�l��]�&p:�2�i"�`�#���._ %��$�}G��$9�q�wAy���u��T�2���>|�DKCp�U�{��5�f��KO�ڈ�
����Hc�`}�;�ru<ޣ�g��v�;$$�7{ y$��A*�ޥcq|��uPR�l��=q�С%��,��pz'F�f6oI7l���G���*M^y#	����ŏN����/�9$�8�-���Z����5��G}�4=Ԭ�[�o�qo���f �-C�?/tI������q�����|<2�ǔ«!N,L/��x������cƖ��������,hb�d�?rUk@���^ rW�C��(c%1��V�*O���zx`��U�.��34o���M ��9` ���[t�vA��X�uy�"#��&��0z~� �&&&�1�=�� km�8�#`Dox���u�{C0U�Jð�Icu���Z�����v��[��92�~֔�x�F�[r�*q�,<��-��	Zz�r\;c��?|)A���-���t%F���r��W6~��W��D7���t�,�'�qǜM)}�u��)Y �z/P��v����\�.�@�u�MZ���9橞�d�r�~�ܤc+uϦU��	�������[IrC�������=����hw�\��_entj"J,!����U�Z�	��*�"K��4Q�4S����
�c�W�
���A	�/-"�!��"1�i]��5�\��h�ϻ�mC�뚥�e�q�mlZ�QZ�5U����Ss¶�����O_ ��]Z���ݩy�5�(�x+DN�#!X�ƪ��7]�^�����W/�J��+2��-6���˷whh����*�#���z��+�B$���;`̱�%R� ӑ'B�bmN㼞�����ih�˺��<�fP4�����M�;��
���A�?���f�%�D��#�"�����	�3 Lԙk��K������Ca��a��;i?�Z�$[�EdT�w�{���C���Sj?�.�j ��fB�����	���Q]mM��k���eaM���]@?�9;��q,�����R�= �u�#\eIO��7fgu �+��FЎ�?>�ϲ���NOK-�ҵg:t�o#�a���d�f�};�<^)��'i��Zn�!cma7��n&���KC������U�{փ�oxΠ��H�|�U�]zwO6��]�����%��s\��z�J���۳��0xď���	�����ަ=�RC��@.�Y�ibb2�=Dg�;� |����Z�5Li*��ڔ��I��֯&�Sn�8cC�eh����c���Kᙤ�f�ɒ���?�����&���K���C���`@^��*<�4d5�!��L��ܢ[�Kj�s:w��W�ܝɇ56����������ռ��"9�r�$s^��s����f�~j�q����
	��4���0+���b�-4]�����/��$v�J>oY�!��@��e{�C�q�p�������g���)���Zڒ[n�E6���L��_�5M�u<6xc*Ʒ6�g����:�58--0-�Ub��^š�R7��"�㌗��G����Ɩ��i����K��.͹�x
SM��C�I4X�g�)��ɬ��7nv宒w)���L�6X-믎��IvD�,/�5Dw���TR�k�yD�ʘ�O5��픷k����Z�0dw�4��8*wFe��.#��o���Bu�L������RI�2y����{��Vk�P�6�����0~���_^v�IT�v�3���Ů�7��<ؼv:r�#�g��b���q�N0�3����#��f�z�syv�y'�h+<�,�SG,����/�tq�����˵�fU�<ciU����0�+ �|������,#-��;���9r�t��#��*@Шn*q���
���zĈ�=rK�(��V�+�(/�����v%g �����7y/Z�����M���r�.�G~Nڱxx�����E?&s��_��z9w�r��@�Kh#>>&�D���M"1�X�n�^���h�A"���pQapo# ��} �vu(V�k���wv
����O*5CXgX�����w�I�j^�5(�"6\tq�`2��o�/]駌��rj���$��w�ET�Q��u����ٱ^Uٞ h��&��7]N
���x�����0�-�+9��,շ��f���`��Ku�b��"_`v������1�
3�? �e��@���8B��P8��(EB^�-+��#:x�:ٞ0�}`��oU�ǉsVC���۪++����>L.,Ց������f|h��;���Ju��LJ�p;طN1��d��Ln��Ƶ_�v�c��@<���11�p�7Xݑ���_�Å��׉6���$o�mK����o0��XR�Wq�;��umY�x�%���L�9�����X��r�A-��|}i&
{�P~Jh%�z8�!�q���!����D׶�c�^k�mi� v6TV�B�����cX�'</�t�y��\w�mu�"2��2~I�r����� ���C8�J^��1�p�2t�Q;qMS �|��u�:$:�3���pSY,u�܋�>��L�i֣ȝ	jj���9�C,��_BBB��v���K��'��{�v������J4t7�ӟ��{��)b��)��#�� E��[�t�`�ՋՄ�.[VJTн��"D������S��?�n��ƣw�C���/��X��J�T�t�[�d���l�� і��^+ypƋ����s�AC����=l^|*��P؝�l����F�LF  �Z�)n�"<y�3�ۂx޺��zB�ڣgjb��sF��I��~��徱f���-����m��I�f�KS���Q�yt����:�Y��Đ����_�S�J/�������жO~�m�D���,�;�L��U��9�D���8�Gi���G�$b�w��#[��65��4�Yex�"������lI����
3��(������+9%�v��
��Uon�1{a�M�'3z�쒷u��'Ak�i<��c��Ќ���>(�!����:��ǟ���(z�*xa||���4�g���\�����:D<v�$��:����PF�(d�
�����&�u��U���ӵ�5{����[l�o�ĵ�le�i������9�M��y����g�ɟܓ��sIwQ�t��4� H��Xj^/a��f�A>��z��V{qhyia����{�Ɋ��P�栰���ٮ�U\®����a	��~��d����'��R�υG�m۶@�� o[��	<�)�6p^)&�/�8i��Ka�!�Z3��$�O2�Ļ`O0*

�p��:�����\��,m�G�yn��y6�3����Ej����-Iy�%��#�pFϥ��03�b˚څȢR.�b�=C���^����
2��D�.�m+������
�n*R�����
�b.�uu�����%�p�X���3�������`CS{ǋ{�6���~1��ӱ�b�r�Z��$���^�1�����b�J4�S�&� �h�*����SI�'�מI-��U5�,c�߹�mר �����P'�8�Gq<A����m0��1ƭ!&c&4r���(�ͧ�C�qX���(������!�����ab�h
����xd�*�3����d�`q��}���b38�$}�&�L[w䅩*�}�0�.�3�'�*�_�b�b���c��7b��9��H��}���^h�@�a�2Ĥռ�Q��I'!�d�N�{�K�/��2�"}�U�D-W�N<�{J��O�=Eyܡ���<eB�uhI�mA�0y�:����ߛ[�V��|�@+s��z��[��"j�"rD�p��e�/����ix��+�-����	����)}{q�?� OSST�1���0�4�'����\l��R��Jg�z��j"�0��˵��B�c���f:�Z�8]Q��\M�왝]ߪU@�6��(.�OVWS%��S��Qg��J��?�m�ݚ�f�/ҟW�=�罌��=l����:X�����ve���j�!2���|�&n��C�i��3 �#�w�:p�?����(.�p9&r���=J��	���2�������m	�0!��˱���{�2!��C���+G��(�e��M��N����N	�7?�h�s<gY[���F�80�&�B�;��~Z=$=GAY#�î_��/#J�R��o��[�,��+�u�]m/q�c
���%ݶ{��s"���ډ�Վ����]<Vi�SU�o/ �U����q�ni"��*��ǌ�j�Ζ�o>�Ù�E-�����v�����/_���8�s���+��? (AۮG��&|d�$�H&'KP�L�G�1ׅS�Ґ@%���b���P���:3Y:Q���`jf��>(��Y�Ϛ:�%)��

��B?!�)��[ �)��k�!T�^{���i,z��7�1�����*�X��v��.�a�:��==�:��튣�3CM�K�6ѭ7��ѕ���c���[:=6t^ii,�V �\F/`P����]�q�v�A�8�Omy�ޟ*���g�n�r{{{��2D��;wdR�-��G3M~�[��I��ן0R�xH��^����,z�}Wo�Y�X4�h�o�4]�W�x�3��d�xP-����z�c������*~�X���0L\9���d���q�Մ�K��`U�̍!୭����Hc/q��B�(��8�Wr�������������D�1����hǃo����H�L�t�l�a��G`5��ngˬ���-@a벦�R����������j��$�k���w߾�Cd��x�Ӻ�C�����h��G(}��ޝ��R����:� P��v�B���v��)}�q����ݾ��zy�����%��j�u���9>c/��J}vS���G���{�dr�Ԁ���x��M�BZ-���V�J�/���jB^��ʁd�ŴD�^�b^�I�����j��g�RB3�s=�5�#�fya%����aR��M���\�&-��������?�<r�R?!(t�Bw�#uO�Y���K� M���&�Ů1�fVS޳,�J����ޖ� ����8`fN�=�� : -׆n�/ �y���?��(�(���_���{t� ��;�^�b�<	�x��!�$��,��TF�튧��������B� �^��Ԝ�;3����� �!�d��2ģ��㪼�"�?�H��}x}]d�Gy��Y�I��\m�H�@a�u娈�u6�|bf����M�n[�x�#�҂�!�I�6נ�9 �0�n�,!�yJ�\5�N��`E�0��WL��ů�G@4��F���k��E��̿j�VaGH6�7�b_.^P���k�w�<�n���{h��o4�%%�r��ʑ��%D�sV��2�8�X�!Z���IP'�n�+C�Hs�e���"X+=��S�� d0�M%����7����[H�����H�;Q��3V��������]���~az�,�0y^.;���F+?�r�i���i�|��\��Y;�P�H���-/�R��@�z0&zsZx������|�n5�20|.�����ʗ����TM�����_Z��z�A7iK���{�6���ߴ�#B�ȼ��m�_�rō$��U&?�M��	��֖t�|��R>D�=��u8��4��>Ы��6��I�Wӂ:��/���o��qx�_�Vh�\�V!�L�yU��K�$9��
�5��_��q���B_�Z������[3$�?~��$/_���Ro��Й��I���.���������)��Fȯu�+�=Z�7�C��*s�~wh�ވc�,rcFF��-:V��ϰ���>O�~ᩔ��a:��5zz� ��/�]OY��z3�h˒���㏑��_Ss��	!B�S�s�-ܩOU���o������5�=���{������N��|�O-�������
l E����
(Nj��~���6cc��=L����43=ʱu�֍B(�?�π�'�Lz@V8c�^8�/_m�������5A> ��g}�Ȳ�
�j��eE85��aM��=�Q��݀���� ����-�4�H׻��|,B����m$�o�H��)�s%��G��U�� �+�kJ���:褷3�矿��Q�Ǒ?~x��:����)}.�c牋nxp���N�@�ͨh�a�o�Tÿx,�7�>���7��� ěo˵��E�/���Evvv���=�^�JއE��!`��|k'�X� v�%jA���S���P�AC��3�e��x�Y���d�Bj�o�N����;e����T���r�������V�Ic�`/�d����ݖ��P�.���)~�]W\^��ۆWq�a����ĉ��c�C��9�n�-H���Tg\�Uޠ;n+<�_8V�ጋ�g ��_0���?�dvV��[�@R6.��z(�*�x�u��2�`����_ӆZ��o���;�J�gb�A�*����y�w�gu��n�}�.s����[��T�.�җm�Ջm�/f�'�ʑ�D#������>DD
.��X�K*�H��g�b��bl��1#I���R�0S�O\^s�eH�~SSSƸc^��^��8W�Ԅq�y'E$o�Hi;�/J�y}}H-O�d���Y����8JuIls��� �f������������}#���E��6�����D�����K������2V�dj����{~�>���_(�kJsraiE�rkeu�O����%��L%�:�H�5�j �O�y�������ru���q���p�.I��I5ndl,ѣ8���0�ή�f5D~G�x��6\,��3�ƏXk5q�m���an|qS��z;�2V�è�u�c�D�)�Ü����8�:K��[!?vg� ����\�ę�P3X������@�q��<�˨=^ ��I�;ɔZ��W=�⮆v�ƚ���{M9�O�~ ����N�x�.���$Dp�A:��#1[=���8����Y̾O���
�\I`�g�D_@�WLb��8����/�&WK[{���46��Џ�]^tz'P��L�K�]�T�C�W�3M	Z��;؂�&?�����4���+\������r^ԟ̛�tY\R^ �"��d|w������ơ�{_F5iuz���E���'�\�n2�8�"������ �b��<�\/�����j=�a=��XLb�^d�-fs}ƺ��$�a}z���Q�[ǟ�V�jx�E$�s[�Bd;�����I�REւ����d�������� �ݺ:vN[�oo�Pd���)�������XP�u��ˌ����D���7�����|��öm�d� -vB4K�d�X�����w%�7_�vK��|��Wg.JV��K�r�0�,..J �K<�j�JIި��>񓓁�"t�/�UD�ڢ�4�q���N�tU ��t��}�O2*��#b�8A'�� ��g�poWw���~%�@��k$�B�ڣVu+�{}|�!N���{a}����������ܚf�d����K���z{���#�S�^/��.�	r���Q����?H�� 
�
k�4+V��]��R�]!k�w��������>�n�x���
��R�q����^��L������[���F���c]Y�H���͗#�#��� 9@=W�K-����?�J���:c� �햞��K��4�����li��q��D�̸�f�C�ALTԘ��s`�G�#`BF��;���{ʼ�{�+ ���]�1l�����А�m��B⻂Or��$���k�ׄ��jP�Z;$�*��������c�Tg�7�-8�{RqT�ƕ�����u���忓i�߮��BV݀$G(挞��ZP逨�-��g ��ݺg_����l2N���i�u_�T��$)f���d��ꙿ	B�R�#����^��C����Kc�_6�7Or�>�O��F�iꇄ�C�Õ�ǗS�ňDVÕ����f�	���V�\���"��L9�)�s�2d��Ц{����ԛD��~�x�|���"�n�*o ��y�GS|���w�X@��͇��vNr�7����It��8��z��U����7�u��ߡ��4}�h���ć$��������m2dҒ4�{�F��3��i�����^��WU"��(w�f�{i�D��a%�;�>��i������5��H�!�+������R J>��uq�_W!$���}�/�G���H�g�����bN��@��-��`�S��4_E6;|�(Ib\=����g�'O� y#��,O��ΑH���� z_feM;�{p�����={���0Wr�7<��A���᯸�����Ĝ�U���DU㪧����pE���Sw�Cpsr8}��(.�s�d����p�n��M��c����7)��C%�.t��{ā�p�S���G��6�)���A?*
W^���,Ǖ�����J���!�yB^����V
���;K���2|���	���>=�k��t�W���C�:�y�H[p�9�7?���=�T%�m�����2�u�K޵W;H��*���d�����[\+�Y����p��Ntv���HL�CC��Oh���_�L3�]6qq��&��ؘ���Rv�-�$9X5휧S���I �J�(O���"�Ms��ϲ��NLL�B�ny�3!�nSn����?��Y�[����� ҆�f��:�:Vc3vK���y"��=]���������x/-#V�;B~�J\����f�%AA"���A�dO�89���X'͑Qq���{�2B ��o>ѦK���YE� ��P	��ςX��E`��׳վ�\������{Z���
�WPs��!q��ﭓ�F��g�tT��q�8��塗�L��02ח��)I����P���TˬO��V�5m�]:ӕ�.�$=�?W^�B�ki!_�(�jJ�5��N]���8w�IbŊ�:0�ZDƯ�Q3s�ڂ���>z��+ql�̰QH�wVQ1����h	%��}ՎZN�����k}��2.K�Y.��k�\� L+�~WI����Yᇳ�v����u���Z��E��A���|9v�>�3��HM�KY7B�Q�����)�UjBg7}7�d�g�OC�7y>�hd�t����l��+���1^�u~S����{Sr���t�*ڹ�����-q���-D$�	��9?�Gx���\���tmIIɮ�۪��g����n������f�e-;S�{j���1[~¦j�ňЎ� �fgm'B�Ta��#�GLT�5{4߀�k�1��2_�x���lpA5�-7E��*!�5���΀��U?��ʉ�nl~2k48L�9[�N�emgM4���æ�B�>!��٢Qv�i���k����Z�-�a�tC:���@;/�C�6�"�V�5�)}sc�L}5t��G��I�������
KW�	˗#O{�N;k���S��>B/��#)�&cUyGSSSCl�;boo{�N�?C}$��H+�4�m�7�n9L�-yYÚ-1�f�5�R+���mA��=
M8�.�_e���V���N�-��{%Bo�Z���������v��`P���w��^���K=�9���6k�h\^4�>֖5��w�?;�סSb�O��o7��l!���,���J�?��Z�[��jJy�W�ݧ�l:�����x'��B���b5��b�Ē�k����A]�y�
�w�qL�N�c���(A$��}��1���hG�6�W]�z�����9J_��7q�jBޜ�@$���@h�ټm�7)�	��z:��ڔ4�q
�šU�*8\{��o��0mr�9�(ڃ���,�x7UCV�{�� 6L4ڂ�pa�ٻ����ރ�P�.�8�1�?p�\`�*��a��s���"�G�kfjۍ�e4�ߢ�;o���.�̷�^p���9���`m�w��\���|�=f�ēi�޻nE�|�G���7�?��hA���u咠���	$U�$Yݰ��$h] �e(��QNe��l ���rq��3g�>-8N&n�i,̌T#��|����1�ݘ��8���_��C� |\	�4��M�������:�X�4dܚ5�����s8��LksP�tlM���wĉ���s7�_��<�1Ϲ"Fp���xM����k)�FXe4Л��	�5��{�-_���d��ҡC��"d���8�OEaJ�27Z�<�[�I	����G�0#��oj�\��$��LOmj���v ���EL蠉V �1ڀf֬vӲH�/@����U&g�>�����So�-r_7<�P���CZV�1U`^��O��ǬL�(�.�Ro?]%H��-K:�2�/��|R-�1���<d2��v��9C@�M�>W��"��$t�M^ֆ�kE'�]�������?*Mj\���`l���(*	~l9�����gC����N"��9��jy#v���W�P�DԆ]��p�����>_��;�����$��K�	?��I�;���M��� i��=[N��])Q�� D�)o_m�=V��	HV	LJ�A�F��(-:j��__�����>�s� 3��5�Q���A�o���O�nL���Y�p��cq~�4�-�+M��}�_�Um���ܤ0!�p�HW��B]�� !\^R7~�,t��	g�y��A|�5�[��6K���dz�S��WT+n	9h��;��!�s���M{t(}�c=G�|GBx��n�h#L��J��y���|�����_������R'a��Dr����������u%Z������g��D�9*��>����0jfg*��0���:��D�J�~\�,و8���P> ��_���J�V20����+�|/�^{��9��W�����H�U+��`
�#��X��y���(�	&��Y��Y���X�Ѧ��FZ�]ǥh[�z�	��㽰�gP��@�u������?idE���L�l?=2�\� ���Kl�9�y�bo�Y�D�Dӕǩ�������X{�UG$ژ�'|6S��T�[��<+n�nS[�C�О�ґ�
t�4������k��ٝ����%�mi�?��A˫%�ꮩ��f�Ʒ6~J��5��0B���r9�S�B"A��J�eV�P˕06J�7���V�C/dO*�coq]�)�?`�?0�m���vN�sB�{�k���{5Bt��M������v��joo��AZIA�"���j��7��)� 4������QvQ���Y��=)���?Tݸ<�z���(�� ���(˟��m��� $U��s�"*� �ݪ�}	�X�$hJ�����+�'$�������vA�(;'�;��%���5z|�Y����^���nP症0�;�����B�k��_�_�L�./�ޒ�3�~��0�n���H(�r�#}.z V� FL�,�i�7�U�5W�hu��Ͻ��Rn��r��՞�ű���w��=�,L�����ڀ�J��_/u��h����8*x��9SӅv��q�@��0��_�kl,����<N(2�Wc�^x��M��Ν-->v+�iW��R�pr���Pe�B�3u�i�&��D4�f;W�	��Q����aK��&�3����Y���ꕂ/�U.#�m�z���K��u�\�ѭf�tq� v^��̀_�صN?[8=�,�p�-D� TQ�6��q�����h/a0r:�o���K:=��wޢ�@�Zbg��È�)5�o��B
L�)��O�/�sQq�۸i�Z��8%g�	�ȩ��nyY���B|g�}�ݷ�Z-4i�=��Q�$0h���ұ�h�@��Dr�۪����VWY)(m�8.�>a����{W�{\?S�"Y�`�*C���QQN�j��憒��V7�a;�A��H���,�wfm\7�e�܈c/�7��7緬���@F���\=�Rc٪t�NH�z�dk�Y�L�""�V�k�6{*�.o+��b���x�Ҹt�:���q% 膗�.��C;��i^�8	�w��GK&� Z}|F/���h3���x���k��ѕ�m�du�!���/%⸩�|�*B���(}��7�
���c���:�7�~ӣ#d��d@$=�Hr�p��Ϣ�T.&�l	 .p����Z]a/G�"}�}�H\=���I�V�A���[vl!u���=��cQ� /n&a̶��!N^h ���2b�'��@z!�٩u��N����Hj(o!��|�@p�\�Y*:�w�s�ه�r�O5�e���Bd��֠�l� ��"��a�Mt?x�N�A�
ӎ�~R���ԑ����dK~J5fksK��3��˯ �+V�`�����S�����ϴgo"�)U���Y*�koQ���#!�$��F�O��ᓟ�\~�����ĺ����.%��%Y�O�5N`��0��r(�ң�:�&���'���y!��̠jP�1ݗW�@�B��}�Î�8N���!�_Ȑ���Y��fЗ#)�D"�I�w�O�+�P�p���F$h-�3�����O~~o-ۓ
y*��︯k�' f�������;�*���ի�k��Tm|D;_0zn�kY���d�ɬg�X)���.�=��|�K��)6�nN��֨[��U܏�nDKF���V������<��LIL���~��~-�UK�p�+���5r��F���m�?��r���>��	>[�|H-��M���[��Tw�[9����_���c���]bnY99ޏ�+^��:��+� �	^�yx]�9Lg�s+��>i蚏��ރ��M/��kõ�m��v�P���|���%S���O�8���� ��tyOKIs/����5���'"5������A�8>�'�"c��y���Hcu��6]'�&*����-�}/8=���~��=�a��G>�!���x��+��p1\=K�,vZLH�
˵i�ʙ'U!W4(��wRpP%�A]uֈ﬏U�	k�3Ȧ��G��L�Χ��oAt�TH��}�-��}�k�jt�æ������BDdP��ƶ`8���V	Ll0|٬pc)��0@t�h6� 8׽G��#mJ|{Vf���r�o�J�OB*v�<|t-(+`��0�aY�W�=�-����4����Roo��X'�AZ?j���m�2�M�J��h�m|��3Я7�8���(q�YH����]У|7µ<ΥR�-�~n�[[k<V��^�^�n�d�<��M�=��� �5�l�G'��üp0���ؐ�f�U��Y���R�=�U�Y�R�K��Xu�����b��Ǜ1���T�\}�����g�t�9rO!�#��O�Hw������Gq< �o�B� �������L�Ma��*��ϥVE��l�U�#���Q?��Ԓy$�����Yy=�S�	�kS������ޒ1�f,�R���a�S�}�~Z��A�F��O #� "���
g�V�`J�_�sBv�m�pVk��DZN�ɑ�sb�G��j�_ꓞ��ў�]Z���Hη��!��%eA�����!�Ç:c���2�u#\�Y'PpҘ��=r0��������;��.�z[lK�i�bL<P�5+�H�7W��gTU�)J~"$�6��L��p~v�~�mD�FDI���ް~�^�m��� ͱ|����T�U��QJb���Y@��tް��)�;CQ ^�k<��w��Q*���!'�%��;�"$����Βۛku[�����\�#.n�dɪ�'(ّ� �yp�}��Q0����A)n���O����I�`7' ^���>S �~�qj;�~Nb�\�?��&��S,,���M6��[�KSQ��23�2�jD_��̙IEٴ"�)�Ԝ�"�,]YHXQ�oZ��t-Y-h��F_���@�U���Q1���}���[QA���=�s�=���9o��D,���v6�w�-4	���s�$��;�ޕ;&xdR�����ba0�lw�:X� �X06�ֲ�g��~-k���=�3�4��יć@�35�^�{2`�xU�� ����W(e$��!^N������OGg�)���Th��-e�A�������N��d{<c���2���mͽos����C*�	�����c}��J���a��b�W�V��~8�Ds��f���@3NݺX
�-+]��v�u���t4Lf�M�q�����+�ذ�a�_���������%T�����N�[�:3�A��p�3���)
Mk&ثA�����ъ���l\j�� &�J�s���UhG+��3x���Go�.7T9U��|:[�����`����DJ	Vg� t��5�ܣ�)E���KI��Qk���D�
�%��q+֠!���ؒ��z���������q�Z����̭s�5Ҫϙ&|Gøn3dE�d�򉼩j���lyzd�8�<�p����G����f߀|!~c�-L�_�-�	��0���Y��~V?���?gum�p��j��l��Ɂnb=�e2D�w�{�>"�Jm�.`'p `��]�1�3>��B��2e���C��
�[ <�(���[��&�yf[K=a ��)ĵ����XD�b����n�{�*/ivB^-o�p�znGx�n���(��� ����Jct�������J�<����pÖ� pPS�q����(�3�ʴ]��<� �4r�Q���+��9t�Q��Z*а(�ji��x
<��� �P[na����N��n��x�/Ù_�Y��mj_֡^�=L�"�:�=*-}0ѶE�A�5���v6d�@Q@�iE|x�:�b����G��jJ�&uF]����Â\m�h�#��n=�G�H­E53E�Xk"lN	M��_�n�;�ZD��9߾J�->�OX��w���e�yW����'�D�V-_�b��PK   �>X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   �>X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   �>X�h�F  A  /   images/cb0ca54b-1964-4771-904a-f612fb73280a.pngA��PNG

   IHDR   d   �   �8�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]	l\�y�]ޗ(:���D�uR�]���ZM]'q�&��Z>MѸ��nݢ���h�(5Ңhc;��I��)Ԋ�;�uZ�e�A�(RI��!^����f�����ݷ�%�����������̛�.R�N�>-����|"���F�'?�Q�Q�P�J e������Y����Ν+R�R���f ���CY�R#l 
��栣(�d�䠔�T��P�Q���쓨���S�NY�
0�b�"	D�(KP
��Ԁ,�.U:A"e��6�W����;�υ-M)̄��!���r�R�La��!n�u)�E��G�e�Nu��f� a��~�e/�m�GY+l�C)���|$a��g:�WP.Cy�޾� %��R!�X��Ua��!�D"���;7==�ppp�J�7(lp��	�P2�D�e��m΄��T@����j�?����v��/;;�6++k1��j�p�B�9�4`(-��+�mg^Gi�'�����!��7����P�B~ p@\�����<���,����������v	
�`�8((��By���K&(I�F�ߊ�u"�TXz_cTLDЇ���QW��S�%	sQfARN���!hi�R��w���k��`�@I
 
�RF]X0�0������򾾾�J��q_`2|RQ$��?�/��f���~U֪���ɛ[�5�y}2@I8 #N�&, �,//o%�+HKK�����TH[˽������C�Q�B�9Ch%�{�\	`�AZ5o�@�o����q�Ii�3g�H%��-0���*a�'dLL�����9�R������Fn�D��^�BZ �\x^KQ�0*&��b���dwww柳A�K~�(]��sJ MMM֧�\�ޔ3�d�nڴi+�>��E7� @��P_'� ŧ�E=' -�_�e��KbІj�' �>))B�üٟ����`"UW� ��+�Y~��(���������`D�$(��:�٦4ؔ�s��m�}/��"W���H�$��36���?J�=I l,T��{ɟ�
۷�� �Tfff(0FOS2��� �-������`��@I������7@cIj� �t�*�&ı6� J��H0hDi;�D�Ҁ�a�&.��p�z)xu�ۼhA(Ð�Ϡ����. ލ���죇��!d;i{֡��!%����R:�
����-�)q�pF"��vآ#^������ǌ{4)u�t��e��H %�ˢ�\&�G�A��Z����d1j��h=F�P�6$�=T�hX7U�<L�ざ�1{�l��9 Z�ragnu��4z{�A��{dl�O ���!0N��H����M�)����r�v�3~b:U'	Ƒ+QJ�12��O+�-h��)����(3`?JEd0Ҡ��(��~N+�om�� ���<�8Q6��8U @ F��v&�N�� �����2zO L5pzTg:=�l&�Dd�*�h:Q�kb���j��-�N�d���TW ���l���po�&$v��}�3VC���-���c�AxV�rb*l ���f�#Km�Or���5�y�#��v0<��U�*�m�N�'��R�"1v��d2�G?�y'@�$�ľ��ūJ=R �X��Q�S* F��:�`؏sb����)�W���� ֗�<@RB�����>19�6Dx��z�������Q�j�'«,b2$�?�@��׀�"��P��'!y:�&|��F�Q:<�T��K��]$�� ������G�\��2�Fi��dP� ���Pτ�I�0hJCo�R!c���2MC�c�	0��w��ܹs�>,���˗�[TTt.�{�K�\%(<����͚։#���b_III�b`$"��������Pw�yԓQZZz�2u�����9s�����&��E~[ОN/���HT���YgϞ�&^�:.���z����7�p�OM����*������;�g�dnNN�������q=��f���C����RH�d҄ �tww��LɄqB��>|����� 62�t�۷�#T=`��]�v#%���Ou���Tv����ӄ ����ϥB!AЉ�<r�Ⱥ���c�����-�8q��<��+�k�׬Y�*�U'�R��n����h׮]롮���l����
�����疘#����������X���P\��+�JJ�����U�V�����UIA���ر�؋҉�j�Dܔ�X:P\�ۡ� ���~
	;�����ח�}��o��MJ�E�eECтH0�����ת���@%Y`Hg"c�֭�Am.H0H�
�h� .^���%K��\�f�AW`|jsq*�A�Ҁ,Z���+V�V`(7v˖-�ttt,K50HS�*؋M�W�ޮl��� _�W�:� M9@���!z{{���!�AzT۶m�bkk땩�M��)��ٳg7!
�@Կ����:����������SҔ�`̘1�F�A�5�cj����G��"�Ju0HS�Q\\�VSSc��"y،�S�N1%R����DQJ��,gB���pm�+Um0�R������X��p�ڦ���@B��6����333&�|0�Cpoi��p�|s�������n���P8<<�'/��&ـX�|�dF8�O�����j2�!G�O�!���!D���`P�>���Ո܋�j�>�*���#ZJ �_ �����`^V�s�PF���Ա�)Xǳ�֡���jD�"77���3sp��(�|�]|����J �� �<t�P�{Lb�kڞ����pFv������⥗^��w_\7L8 T��W�S'O��?,��]UVWPP��i|
������r���'%e�ƍ�{��~	�#�r.>�`�'bB2���6m�g���*�3�������ӧ��1�Dn>�\5tp���'�����Z���~��и	� 1@^~�eq���t�D��2�����{'9�F`K!��)�� w�À�}��v'�$�2��@��#\NI�/�[}�E��^��B}����*%�B00�
蝰�SD2tb�Ҡ�+`۵�x�߻)%��b��S@�;�(�{�d�[�6�n|	ݘǿA\����?��},{
Hvvv�5�z��!�6�a�9�"ˠ��u��W^yE�u�]QU�) EEE�����%�ħ��A<���ܗ����3�׃�ak���s�Ԉ��x*��Ə{���ȵ`QW� t� ~�c�S��;�ݬ@��]�������`!~�ɍ�s�C�Z�	�IM!�m&m�9�D)mg��A}=Ѷ�3@�2`v6DFtqqsNN��`U��r{
k�������p�

��nK-��]j�	ڕ�X���J���y�e��8��n�v�W[[{�}�ܠƗ̇dT�*++���'r��\�s��JrqG�X�Z�r��>6௮�N�w�[9;��?�ݗ7�f�D�ZE�w�	rcL� Q��3@`�Ekk+|Y�F��������=��Q�� �8��uww�#��]W�)�t�j�c_���,..�_Q��i �iН=S=R' `8gA������?%rY�R���(AHI�ta��k	���� ��%��\�pNC�ma������%j�J���7�|^2�F�1~�����|	'n�b�����KP T���+w��2��+�3އ��+��#��P�����w���:�NL1W���t��"�|�^6-:{�,Wd�1����ӧ��+`�4�Ch�BF����"� ��\���G!L����l�(ޅx�G�2כ/���p�677gp�u��f̰.e��,U"&���Ioii)I䫁"6 N�"ҲS�:�u���!��h�P� �/;��C!Eڒ�dS�����`�w���b9mkW�Ĺs�Z�W(G e�	��C�����)���-�����xYYY�+k�
�O��h)!��!\iB}ʆ���q��:TU�(� D�AG�����FK��p���%%%�)��ȕ�#_�4٤E�?��������[�pa@�G�l'��9�[�lY������Z>Jܳg��3v���+�.�:T_g���5��KOO�80�@���a����#q���6�F|޼y|gT�����������j1s�L���'�M���lc	��ɷ`/^��H0(8�'���ӽ�1��V��Q}=zTvl���V�8��QGP��SlE#7}���TQN��g$���P��s8��P�Z�*�x���a#KKK�r�������5���JUV�	w���yZ���}qD0��MqX,� 8�k��>-X� ���L
���!�>�G���*P���:�w�^��c�´4�����܉Ɵ;�Lc�M�^$iN>h�l�'��?�s�Μ9�O	vzRtH��<z��!!�7y؉�_��+W���M� d�Nv���.�@ 0���lV^^nƎC�1�Q��j�Imܔ��+U敽����ol`.j&�s9O&�����Q��ީ�N��`(�
;$r��X�U,+Mt�fԎ�,��!JԙF! �+����DG谟#T�s�q� &	-���rb:SU&Y��z��ĲzH���}0H8o_Ku鳉�ca�y_�LZ��S/�r<4J 8��B�z^K�/_�N.Rd���_�7J�dHMM�%��N�q����������3��t)/��u��VF�M#* �-}�b#U�M���7N3U��
tvv�.�	DEE���@�X?�Ƴ���J��X�"nz��-�Do���>����2��%K�9�#2@�ljjb�����f�� (d�Rj�˵�K���)|ǭj��)=A+x�4�  ����H�=0A�A��p��=���</O�� 
�N��ןm\�f�ZF�A���F���1J9���||�ɓ'-L���[ޙ
,y��A}���.MT{�^�S�Jq�:�������WI`�g��|�P����ӳf�=N��<UY���v��|���:�`0A{sJ2��5�L�����Ĭ MT)1��g��ըU.�ܓק�7���) �3�K�:7�z������	��G��=��hԾ���Y�ٹݻw[^�ڵk-�n�)���8.�P�%�HWF^3�]�0��|T��|��S3}&�;�cǎ���F���4~za3���>-&p�֦M�,�N�F3R�G�D�p$:S.\�$B�,�$1T���ie(��4�6�^RR6�$#�:c"��@���S�Ȯ��OR���؉��� ��&�9��;Y��$s'KZhP?��+��t��~Ω�ɶp:ٓ'D�A�8g`�D	%C��Mi<Dُp��a$�m۶�֭�s߾}�p�6�������^��5�F7ʧ(o"p�T�|�����G��m���i��$S`l�^|�E2�=0`�jx3w�Ӻ��.���� _�}���O� PJQ�;0ο��ߢ�?���/\��o�P"1�?w�Xr+
nIэ�C��YpO�g I7U�CxLzL#`ހ��Dk�K��x�[wL��h~���;<�͌x����~�j�G}��<DSW���Z�K���ׯ_?�]|W��H�6��IJ�Șb�7�x�/�S���xb�������:R-V�5��U��|��	���mo�t
�^�-� ٰa��N��K��hW���BOS��!�C۷o?B �9d�Ν;9s���Uu���=d�n�&�������x	J"�M��;�K��mLCu&�� 	TS,,�z5�@���ǤeY��~�l��*��Q�N��!y�ózF�/�w�M�qUA����#�Wop=�Q�\%��_�\_.��x%%q� �N��4���0�P���;���3A����(;Be�^[C0�m�_�?��m�ߠ���/(q� �P�����E��k�?!K���wI�ek��;��Ư��P���xA��(?G���h�)�#D�M^;�;aK@8��Sn��^��h�b��ⶐ�}~]�eyh� 0h�~)�����fV�����r�N�1<�.�\�R�r6w�i(O܋}'�(l� fP��ghh k/����#D�9���a/2���0�i��Ly���ۤ��i�?AYcp?��-y���g,�DH0�)�F�\ AC���_6�����BuVch�<w�K}_ $�r��l�G�L��d�1�b�����u�Z�b��?l}j%=�?2��Ca�7��B5�D��3�<#�x�	������-۾Q������Ai�h@1���h$���(/�z㴀�{LUԵ)����o��C�O&n��;T׏���=!q�*PN�)(�����h�����G�F��+&��������"�)u����6�A(�(l�}�0#��nQHJD@`� �%����^�e�\�hP�dP�~�ԱGyD��M^�5�z9�Y���t�ե=)5l+��"�nR�v%, 0Jeū�9qt�.��Q|��p�`^�dA�"z�5n���m��d�c�=���S�t�ɋ/�������JH@`p%;e��)bҐL�V\D�&�>���{"zzW^�KJ�m��O���~�m��m ��CJ�5��qLp�ѹ��Ы�9�+�N��������3�֧3�v��%l�����Yؠ�j��uy��e�8@40�8�]�����
��-�@8�i��f��/E��k� Y#�r,��u�B���S�J^�"lUr��@��(�
s�'l�oV}oξ幜C��k;m�-���ʗm9�"(xTC������p�?
���P��8�7ܐn28�j0lt���%�C�Y���g��5 t��8�}�����C%]Ј��aN
�&���D�0�O����I5L)q�j�&׭�< �<�A�c�a~�Eqq��5u٨��:©�
��l�A�'�s*�ݦ&A\PhS6�)hI��=�4��\�C:(B�����%]mp��L�H\�'w�`��r�۴ô~(T����A�2��m!Ϲ(ĪG��o{%�	�ø�ް�2�;�{<��C�a�8Ki�s���
�쯢�/�Vސ�	���Q@o|���̴���]���@̰����wĺnw9�m����T� �s�\˕w9����{�+@����$SѣL�c��3�&����ã�ئ�B�~Sr��W��,܉�g��$]^hB?�!m@��쳣��"a��h��z/E��^�Ʒ,�鹲mGb��s�B�F�;�r��G�za��3��7����i����^.D�u���Ƕ��M����C	���z�D�ɓ�t�E���U,08�db��:ݖUxx?&69��s�����ɢhfo_S?�QZ���9&�'�:M��RB��̹��% ��Cu#��d3�3�{2�ӓ�"5P8
�C7@�'�?�S��)��{�H��s&�N2i[�d�t�@�%1wo�mx����ݲ�R�P���|�I5ZM���lw5MJ��=���~�U'��v_"#2�c�_p�\� )F�H"�~3�$���u���v    IEND�B`�PK   �>XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   �>X�1��8  �     jsons/user_defined.json��n�8�_�Нi�W��s�(�&m�fSEQ�0���AQ��e��Jr��v&��x�X���9���?6&�Meʯ���¤�4�n�*���3<#�R5I۵
�_~��8S���E�6ya'��Ρ�V�������ui�-�ҮV����@��8�L�*3r�P�&�c��I�5R�&(J�H!9�;KS�2�Խ�]��\�u�ia�"�e�xJb�T")Mh4�B+9���\�-i	����^Λ�M^�-2�E�^��f�~������tٵ_�ۮ�������oӏu��p0�m[��w�
ZxJp{#����%<�벁�Y�Ĵ�>�}��j�MǱd�������=�x�ډ�C���^���N,bC/,��K'��ҋ*�L1dF^�7g�����b/�%����J���d�C���L�^�C[Q����n��T�o�/�:��[��E���B��C?�1�R�$���S7u�Q��\��#�"~�š $C[��=dV24a~�%9����"��6ٴ�/�mZ:�i��Xw�БMKzbc7udϊ<���:�X��>T�=F�'5tS��6�;e�Ⱦ�<��@�#����EG�.�Iu����]�'�m.6�yIO*x�;�~�k�ۼ���<G����C�Q�#�gQ�%pvO2��N˶�Mi7���m鰭7�^(���b�)ڲC���� �8l�[�=������]o����e^���ܷ��[�������FTE�)]7%&���g�P�#�0E}���"0�kumN-�I}񲂟��Z��}������|��6��V��O��`8ː�T���Ri(Q�	&F��Qx�y��KSF4�ƱF<��	!(K���0F���7M��OO�CU������2kW ���?�2E��hLf��]yx���/3�7���9XG����h�j�>ֶ���&:���h����4�xr�ظ(�#����̹�t5��Pn�T�|&h�e��~W�w��Y@}89�.ޜ�x��b�$ՇO��2����ϓV�=�Z	� ��Rc�P�%���m~<C�]�*�j[�%̉�@��6�$�$"D�Ran$B	d�8�:�B�ƣ
��P���I���JB&��)fq�E������ݚc*�Q1��@����#ؼ�<�dϮ ���tԠ����ڦ��~��B��;��s��sE?o��=�����ǿ�l���-S���b7�'�2��q�.l��Z��Ѯ	�H����~��O�_�}Ĺΐ�9k։)'���Di��$
�S1��z�ӱ�S��i|)�&R�1A��<��c"��D8&�1��pL�gM����PK
   �>X�
7 �  /                  cirkitFile.jsonPK
   �>Xd��  �   /             �  images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   �>X�]��N � /             �>  images/907530ff-a8af-4c9a-ad67-f4101e76dea0.pngPK
   �>X	��#u } /             3� images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   �>X$7h�!  �!  /             � images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   �>X�h�F  A  /             �% images/cb0ca54b-1964-4771-904a-f612fb73280a.pngPK
   �>XP��/�  ǽ  /             yD images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   �>X�1��8  �               �� jsons/user_defined.jsonPK      �  8�   