PK   �?Xu�ŋ  s#    cirkitFile.json՝]o�X�E��@�j��C���5��CwP���$ d���XY�TM!���!�X���Y��J,��K[WG�$�Lv�_ۛf�ݵͯ��v���\X}6y�ܭ?.Mg���f�m~�-?��\��?O��h���v����}��|1[�����rZ)?;/Χ��Զ��)�R٤&M.^�={���Rca��Bj�0CT!5e�!���*�UHMf�*�ff�*�ff�*�ff�*��<�U�5*^(��(��Zi�b���r�����������������������V����������f�v^�>l?���n��~�@�a{��m���o'�W��E�����?loڛ}�X��*-���������y���fW��z������+��𢎼��	��x�/f�Q5{U7�/�W�.)��%a�L�.	Kd��wIX"g��wIX"SĿK��"�]���i�x�/���a�L?Kd��qxX"S�kgX"S�kgX"S�kgX"5U�v�%2E�v�%2E�v�%2E�v�%2p�7^;�x�Kd�x�Kd�x�Kd�x�Kd�x�K����ΰD���ΰD���ΰD���ΰD���ΰD� .��kg��a�L��a�L��a�L��a����3,�)�3,�)�s 1�D[z|�6pޱ�`$~�/��l��0�8]ʂ �#�����bz�}a6|a1�
����(��t�)Y�J�;��X��\X�*�;��X�|��zW�ޡt���cֻ�Jg,]j�ws�;��X��,X��w(��t�9g�;g�C錥�{3��j8��|��]�����|�����p�`���;ya�������� ���I��3������g0����'��`>�c�N,��|~�=��<X>��|� ��>X>��|~|��,��|>3��,��|>�����A_����d��i/�[�� �����;�����g0�O�����g0��YG��x*'��y���//h�~
8��|���0�?8��|���6�?8��|���<�8��|��\B�?8��|��,H�?8��|���M�?�/�&/8��p|)������sfa�������}a��/,��|>O��,��|>���,��|>7��,��|>�������g0��Ǉ����g0�w�����g0��@�����g0�wo�����M��Q������g0�ẁ����g0��������g0�w)�����g0��W�����g0�w�a��������=m`��������x`�������}�`��������`������罛`����dw8�p����������`������睾`�������=�`���������X�fp�`���p�p�`���v�p�`��|#��5�nIl��F�#w?�:�u`l���� ��$G�� �q�ӑ��-��q�ё�w
;����a�&�������:pc�?��;v�����6v����V*{��EkHE�i���:�����?X�k����?X�j����?X�i����?X[i�y���3z���]��U1�ΖE;���j�ȻN������^ت�ʑгv��Ӄ�Y�wc�S��/̽�^ow�'Jݟ��˅���f� �n�n���f� �nAo���f� �n�o���f� �n!p��g� �~�p�DrU�+�X�6�pSJ�r�V�+ޔR��8Ą�o�
8��/C1a5ܰ"N)�K�CLX/�:N)�˗CL��7w ��񢫾?�0au�諯��A&��]�=oSZ�A&��]�������LX/�:N)��CLX/�:N)���Cq��%V�)�~!q��;�J��x��SJ���V�K�x�R�#���:^bu�R�*���:^au�R�1���:^au�R�8���s��Iq��WX�����!&��WX�����!&��WX���EԡK?X��:N)��CLX��:N)���CL��M��&V�k��SJ�2�V�k��SJ��V�gX�����!&��ϰ:~J)|�����C��=��p5w\c�펫޳ώ�w@�:\��q�x��
�W�pEwƁ�Y�*諂u��;���ls\�U�:\	�q�x:�
��`��8p<;W}U�W�g8������*X���3�f�UA_�Õ��g�㪠�
�����"�<�F=t��\�'��eIoE�K����󲤷��%�}b�{^��V�$�i��</Kz��`�4\���%���0	m.R�˒�j���6��eIo5qLB����󲤷�H&�MÅ�yY�[M,�ЦG�ؓ4�LBk��h�{�[M.�К���\i�]]��b�t���&�=AK˒�jrY��eZ���\>���\&�5mz��=��0�wvHh�)Z�M.+4�LBkZ�#��V��$������o5�LBkZ����1I��$������o5�LBkZ�C��V��$������oEw+�nW��R��JM.�К����k���2	�ih�ǀ�[��2	�ih�W��[M.�К��{>h���2	�ih�w��[M.�К��{pH��4�LBkZ�%��V��$�����(o5�LBkZ���V��$����5oE3�DS�4����J��$�����Ao5�LBkZ�}��V��$����No5�LBkZ�E��V��$�����ZokM.�К��{�i���2	�ih�Ǚ�[M.�К��{�i���2	�ih���[M.�К��{�i�u�����Z��jM.�К��{j���2	�ih�'��[M.�К��{Kj���2	�ih�G��ۙ&�IhMC�>5�jr���4�޳T�&�Ih�y�#�>��v�"��ʉn�c��FT����iv#U�^��4#UNt��r��H��G����<v�A����}+Ì�SK���9��}�3�O�9:V���+{�O[��Q<\�p�T��Q|j�ʱ2�(>��Xf�Zqq�3�O�k8�[��ŧV|��l׫vU̧�e�N����.�´\ͭ^�녭�o�<K�a���Y*���O�L��6��徝\�� ;~9 �ꦽ��ׇ|�W��R�;B	��=D� �ԍ�J�3B	���!��Rw$�AB�K$����AB�K+$���ÔH�jse�ۆnJ)��a�j�aśRJ}�d���mX��R�&��V�)���u�	��V�)�ԟH`���o� ��V�)�ԟ/a��:^`u�RJ���	��V�)�ԟcb��:^`u�RJ��/&�cu���8��}c0&�L
w*��%V�)%��1au���8���$0&���X���Ƅ��
�㔒ϗǘ�:^au�R���wN�;)���
�㔒ϣŘ�:^au�R�y�V�+��SJ>O�����㔒�KØ�:^cu�R�yPwu�������㔒�W���:^cu�R��V�gX���~|�	��3���Ro�`��������$���۠UA_�&aM�`��
��`5	kj��iU�W�IXs��:�B�8�`5	k>��:�>�8�`5	k>F��:�:�8�`5	kj��iU�W�IXS3�3O���*XM��|yZ�U�jV�'X4�KBkZ��Y�(u�b�&w�&x�&yIhMC���k�դ/	�ih��y���&�5�����V��$����9o5ILBkZ����V��$����9%o5�LBkZ���V��$����9>��\&�5��U�x��eZ����+���+b�Kb�\VhrY��eZ���8���\&�5����x��eZ����D���\&�5�ϭ�x��eZ���Q���\&�5��u�x��eZ����]͍I�\&�5��=�x��eZ���j���\&�5���x+�[Qt��&���\Vjr���4�>7_�&�IhMC�=4�jr���4��+A�&�IhMC�=4�jr���4�޻B�&�IhMC�=8$�V�\&�5���x��eZ��zO���\&�5��v�x��eZ��z�����d��d�\VirY��eZ��z� ���\&�5��>�x��eZ��z'���\&�5����x��eZ��zO-���&�IhMC��4�jr���4���L�&�IhMC��4�jr���4��sN�&�IhMC��4ފ�|��|hrY��e�&�IhMC�5�jr���4�ޓQ�&�IhMC�%5�jr���4��#S��L��$����^�o5�LBkZ�Y��V��$��<ڑkh��t;vu{D�D7ٱ��#*':o�T9�+{�ʉ��#UN���r���H�=�ǎ:h�2��Ԣ�ce��{jiձ2�>���Xf�Z&t�3�O-�9V���(>�J�Xf�Zr�3�O��8V�ŧ�5��ˌ�S�>�\��U�*��ٲh�U�^MYaZ��V����V���j��°|��,���ӧ������j{��5��o���l�q�ko���U�n67�v�nw��ׯ�@��������$u�ľBV�������h@���C4�]$�8� Ό{��a�Y�T�_�7b����}�������_s�Yެ��<�3h������M���U�	�齃v�ߍ]���w2�޳�@���CE	�+�]�@���K)�s���6����̟�^]����o���zr�G��y�h"��H]:	R�%R�n�a�ԥ� EX"u猃a�ԝsR�%Rw�:H�H�9� EX"u�̃a�ԝsR�%R�>Z���I�O�~P@����� j�E4���Q��PH����� j��4����?Q��@=�k���S��8%H�z�] K��A,��vԎ�� Pm�tGXu(���#�2�����q��_��r �� jq\#��@�1��%P���%� ����[Ƕq��p ��m��� �i	�Ӹ�w�8�zZ�4��� ��V@=�kx'��8�J�p�i�Ӹ�w#8�zZ�4��]. ��V@=�kx��� POk���5|V>�����q��pW��KX@=��z��� POk���5|&'���PO�>C� ����C��s�Sx	��g�pm���|�[�H����ݱ��gqm�|�����2Y>��R3����!��|��4�7h�|�,��|���o�X'�zY>���Q�ߠyN���|�f�'��C�c��K͠�����̗�A�N��3�����@M�wo��G�FM�w���I&4��=��Lh4���K{H'��hB�[���N%0�ф~�5�!�L`B�	�.q�C:���F�tB�	�&���i�M�3��tN�	�&�Y��tN�	�&������	�S�|}jJL����-0�Ϥ��%[`B�	}��![`B�	wa<���̀z�t�G�SLA���hB�F{H���hB��F{H���hB��G�.B���hB�OH{H���hB�I{H���hB��I{������Eǖ��-%[`B�	}�,�![`B�	}�/�!}�&4���-��9&4���\��9&4�����9&4����VtN�	�&�y���tN�	�&���tN�	�&����tN�	�&�����<|�
�S*:�TtN�	�&����tN�	�&�~ ��tN�	�&�^&��tN�	�&�>,��tN�	�&�2��5�S`B�	���!�S`B�	�w�!�S`B�	���!�S`B�	�g�!�S`B�	���!>��TO甚�)5�S`B�	���!�S`B�	�G�!�S`B�	���!�S`B�	�7���)0�ф�W����)0�ф�����)0�}�p�␃��c���?�G8vE���O,ؒrO,�b�Awӑ������Mt���.�cGWxxF��p��:\nm���W�X��0�L6V :�����0��5u����X�p�����Wc��t���X��8��4V :N��$��>�V���D��zծ��t�,�iU�W�E�wZ��V����V�׎(��������������~���l�o}i���8�x=�����ɿ>����_�|��[��|�p�6�-�75��|c��77��|�nI�nE���=���ߣ�=���ߣ�=
ߣ�=�[��l���o�!w�7��mh�FYnp�t���U����G�og�:w�|�p�#�-�<�>$,��� ��[V�7��hE^^�Q!*R��>�������������s;�{�����OM���*�*�O��O�ç�����S��S����us�77W��zs�wK����l��wwm��l�۫}W y�/���-��,�G��O��v�ߴ����7�����U��w��_�7����?{6�uy}�?��͘����f��&�_���q�Ywrq���m�����u��]��w�]��\�3f������j������� 7; ٭�67[�$�亲�o�ه���ūy}0��lQ����5�֗u�ߑy]��J��2���e�����������N��&��z��Y�B���>�lw����	'w\{�[]�������U}v>˘��T<��8xb~�x}�xu�xq(����~��h�������ã��6�W��jv6[��z�7��Ce?����3�O,�<^<^
_������,��=<:x���o�7�_������f��=�ث�U�u#����/�Nճ��������_?����l��bV.f�y�gqV���|V��y�Y�e�L�M��z>]�j>],��4I.���l��Y��g>糘?e�����=R}��4��iU'6�gW��7��]]��/���l�Y�\�oQΫ��1����o���ͺ��m~'eQ�꿄�&�W��$�<<�q�޿��W��k7���-g��;���G�j��w���/_�?�����nڏ���ʭ��&����ݛ�śɟ~��w}39{���r��is��u�ԋ��;��f��T�����-?�L�f���h?l77����w��o޼���?�~�'~��ĭ?z���?���4����op��V�OoU�K6��h����L>���x�����?T�Щѡ�8��C�����c������s����?�*�d�Y:��O�gT��$dt��o�������4?>�%z4=?v8�����*�=�X;^r� �Q$0 f����P̟3 o��
�,����c�ѧ��ox��7�e��c�So��f��[y����y��Mi�҃�kG���	K�{���ũ��x�Y��a��^�Չ��ks}����-��n��qEy��v?l��]�-������ݷ�o���4��oPK   �?X����H   C   /   images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngC �߉PNG

   IHDR   d   4   |l��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��|yx����=[2�=dOHB6H���Ȧ�
����R��jk{�t���zi۷������R�*b�V@TY!@����=��d��=�L&$di����I~�[���g��9Ϡ�Y�����b�x�Ǉ���'NwC�R�j.�s��u�B��Z�?q�'-jJj��c��c¡�v9�v�w,��G�O{5:L�	}xߋ�mgI34�o��RB��h-��%C����v��:as�q5��Q89O�2{{Z|؟����,{r��
�:6B�U������B̞1}�������N���*�Z��Mya�������\.}2��Á��V��P+ZL�o5M`�����3�)++3(o۾� ={�ɖ�j,tOrL�_�:��E�]�����������S�qy��Mʰ:7�-Σ	��my.�cA�	Ĭ��Q�Oar�e^�3<C��Y�e��w���k�5|���Pw-��X�'V翐�����mGOgZ�.��e����@�� B�@t�Q�֪eR6��f�賸au)}~\���e��^\���RM�����FNz2�:��i'���G���E+�AH �F�9D��59�X��5;e��DJ�V*����8~z�ɷ&'�{%8P�����V6w@�V*���j4t<5!6�ʖ^�4t�	Wx\HU� c�MN����H��BhH04�h��h�Z��׏��v�jơ�N�t�`�0|=0,�H�����c0(*�I�t@���p{!���1==�s�0-k<�b���@Q@���fC���ӭ�8^݂/��Q�a�٥5�"96�/k���7O�}s[��*��,�AV豿��������7�"�X[�������i!��T�wAI㓑7m*V,�A�ށ�GK�i%���p��Ac������D�.h�k�W�I����~�(��f�c�iț<������zss�`�utuu�HI����k���U���� �m���Q�D������*�
n��Wb�j�3�
��	hii��`�
!�������T���a���������CxsW��c��'�e�A�ų"`�*Fŧ�jZpOON�����W"V>/y�%!xx��#8�h)���D{{;��܌��^!:�����0aRRRI�187%%a��|��{��8��.�O��9��zΚ��-�I6���+������������ݻ�u�V�<yR�Ɏ�d�J�PZHFF�.]�U�V!++	I����k�?�8�����e�U�5Rg�w7Y�ƣ��	�"'#���?�>���
M&�yY�F�҅�����~I��r~pЌ#G�࣏>�W_}%��K��S	�������E��zsss1.:wݴy�����wa{�����I�ya0R¼x��B,_�� X�"�oߎW_}� 5�e��F=:G��Y,�8q���X�~=��<��Cb=�����"�����r�Pغ�f^��һ1))ڀK�C����}&|Yg@u�Opc#X��S7��{�,CHX�X;�?�	��n���3�*��+��y}�x���
Q�w�yG@�я~���Lg*��X$��ފGڅ���9���T<YƳ�Q��Y"q�������q�F�8�d�PrK� MVE���dF?i�iP����_��_�w���ϟ�I�&�?P��ڇ�]k�83g-2���Rf���$���g)�C.L�g�ñ�%y�B4�9ߣvS�䖟X���X)q�l6�7���/��Ʉ Zg�&�ؙ��
^/���t�J�`��[��o�>��7��ʕ+����_~�k�-��q6&�&�f���ibFSS~������iub��� L�LG�����F&Ǉ�h���@{[�O���|�V�Eyy9x����X�b2H{��ף�孨��H�c0��`4ۄy�"#)
��:8u�A+ٍ͋9�0c�x�t�CK|>6"�m��n��¼t4wP\݊�-2�G�����߂x�n�Y8��r��100�g�y���D��`�൦f�#�,��(��C`��Bz��q���vY�^�Ǐ�cqs=� b���Խˡ7��%6ӛ
�(f\+��������i30uz��G1�?%��9-@�]\,�f��T)�ع��� �F#�q����Ǵi����v<��ð�Ւf���z�"��ff�AO���!� ���us�VbޔT��eAv2��}�
'cJZJj�x`�l�,vܺx�\s��E��?�Q���o]���q��>��h7��C��&�!o�L�Q�~v��1�x ���D\�R���܂S�J`"p���{N�����GJ�<~�BԾ����HLF��G*��U� <"2;v/~0xL��M$���?�ȄU�O9����Y�/Qdm�������(!�_�BX���������n�K�Y�y�t2o/lD���l�l[��SR����퇫�EI
rRĪq�dQZa0�SSq����Z�;<XK�ha�9d^��5��ƙ4�	���� Afdgaz�,YӅT�����dM�QQ(:p]�bM,K&9�/F��<ܽ��o�aG|�y�z�Ǎ��fbJN���mۆM�6[��=u
M�-�����u ��i���iBPp%N��I#<����7^}�>�P��^HB(������=�P0W�jw���G���0g��N
�UL{�	�����ാs&���6��d塺@Y���:|t����Š�!�E����)QX4o�ģS�Nᥗ^b�H����s|5�`��
�u�'H�3���%2��x!����=��)S� �<����`��F�u��s�a@8�'�����>�'6,(�C�I���IS'K��+X�J�H۬V�\32�
$���<AC~ۋd���q;�|��K��c�	|7�p�fcav�QL�B};�,Y�6�-���pk5h�6�bs�����(�m��RJ�0�,�&�<��M[(����u�`�,C���f�x1��^{}}}$�-��ř��ȝn�:���!�ޡШ��{Y�V���B��OwJLe��Ĉ�����3SQ�I�0À���ɈFf��{׮]�Y[8�O�1]bSvO+�&8�%��vv��7�L>�4-��$��T,�����g���Ѽ6��P޲���֓� ���LEc��fsbDPf+9R�$����Ҙ���51|o߀e�^!I:̜�-��4~�Ν�r)S��|!*~ː�@8]kHl!�TС$r��x�?b\$&Q��x�����vYI�����{��c�Q}���B�<2����l��ux|�NԖՊ���\��`�X�� �W�J@#Ka��Қ3o.N/����~]]�$Ry�iH
/BC����$^�)J���tW94'���G�+Z׬�����?���az�������n��p�.X��;�e����jQ���Z	�LKANB�֛I�J l�Q:%rғ��B�؟2�<A~�
[�m�B�g���_�j����3y���db$��u��=zT ���AV\��p�5��C�ʃ܌DZ_ �/��R\1��#צ䎥�u1��3� �:>�aוH�My�S�$�˗/��w���}>�bB4�����\��:O��:�؂�'Iʔ��-�27���ޞ^�EF�ű��H21���Zy?+ ��MYc�WjpHP"5!F��K�O�<)w`e.���\�^��5)\^���K�Gme����Sl���'FQ���k��R�@}ȣ��U\	�I����Sc�p�e�����5(�
����v��V�K<A.Nr�NK~;n\���Tx�еJD���ߜk��b�j��Q��� W
�m���?}����}��a �{�A�/TK=����%�`���ݗ��QA���6��5�`.E(����X	t�@J��[׉����!-�r�w�}�af5�!����u��Ā��:8V���rrhw�`YBۆ�����-�@��O�Juق��:���pY��D����|_�0z� p9}�Kz��{����0 V
B,,h�����5ea-%��;i�<h|��XK�W�9�:����؛�{����8씧8�\���������/!��'��i�)��}���X9q1��N�P_�jw�)��Ff�qXOLL���o0צ���M�R��C��;)	�Sk~'�D�tW��p|%��D����c6L}�UV�v��a�U�*�4�r��^�N�db�M.ޚ-�=Oo�	z>��D��ϻMNt�(�NEzz:"�]q,��%ם8��=�)����b�F��Q¦PKi�=�շ����p�qM�,\��O6�=h�����ڒ(q�0V�F~���+>�
	̸��� ��2q����;?��w�."8��}p�)��B��Yݨi�cf�4����P6�EEF���q��#�&�G�'�����)��mX`���K��]�b���={�\�Mϭ�0�J��݃�is)P~�+Ic�����L���66 ��U��O%�����
�`W�J����A��FC*�{x����%��l�����cٲeؿ��.q.\ ~����,#-3�Cp�|��٘��.�x�:�a�:�;l�-s� ;;��@Em#�\���"�c�� &6Nji����F�]u8y	�q|��[Ɍ�uaP���rD��$���5��g���Ȁ�hjmC��$uAëf����Pd�p����E*��z=v~�V�^��d)D�R3ӥc&�+Ŷ��S���N>��gS���r
g����K��j1c��Z��\Y<�&V�6���:,��EAA�Ν+JȊT^r
�/
���J�Z��ű�<W9X�آ��J��bs��Sb�L�V�^����1v��
mnz�Y�E��6�����Id��3�>� ~��_I�ݻ{�⑛7��Cu����}Z#�`4�IBg�Х�D����<!+e��Ipsб`��N���{�;G5�.u\l�$nڦ�����;3O�G��?���Ue����c�C�x).(�P�������ix,�_�B+[���>�2��6l/��-QC���C��6��wO#3+w�y����U�-��$�͞�#����W��9Fh�>6�4�Y��Ox���C�슷�<���B���Al�u�F�9E�1�s=�� V�E�z��'۱�D��?Gv��{��K�PY�I!.ܐ��s"t.~��G^/ˢ��hnh����~&ۣ�7>���hTg��(��M��N6l;���(�췿���5������o���� �����~�Q�P=�'�A���ȧ)~�q�z֬Y"ރG����U4g��gh���k��i�F������T7wK�W��C���h7+�����JCTL,�|�I���ٳG@9q�X����dS��!~|p:QT���&���>�(n��f�7����]�{U���O� ��=Ԅ�̃X{�R��*6皚i��۵ՕU�6#_�V���=C�Tu�:�(^�46����@��׿���.�����K���::v�ă�CT��6�GZ�	Q����'���'�s��[��C� k�	ύ[�g��rf|�?�{�R���?����,�RGk�loGVN��Wt�[T@�(���O���N6=�e0�������\<����l�C��<��[������,B\T8
��A^^�~�mq/���İ�(���>��01��p�0P�����8@ԸG,�����yO[�ڵk��v=^ܰ���"�Q�F��I��w
{,r���zS'QgàPU7�E�E�D�t��}=s/2T�%��9<\�4�����<��|V��ؽX�l)�������f�͛7����?�*O�b%u�Q�E����k��$����o�y��`��!�¥eЄ�l܁��]R�:{��e�u��y����4�ysfc�ĉX�n� ��[o�����4�Y1BQFm��I�֬Y�'�xBr�yԞ_�16��WFvC\�	"vc���[G��99�������ơ��$J %%�|�ь� -��c��/�)��{_ɽ7^����b)LO�Cp��˙<����ԐG�[��pn�.�c�op��u?�+;��R��A�%��_�T�O��9�6�K
%���?�Nז-[�^__/%��2È�[/��-K���1�PQQ����������B�������;��/��~�_����za�!.2f��p�NO�����X	yK��y�K���ݶ�Z��p�s�=���k����QUU%���lο^�e����[n�E�8qŃ�b�{}�gX��	6������l�A�����QZ���+"%5E��2[`Z����R<�dq��� צ�<����38�I�~v(�+[�q���ۊ:ƻ���Ĩ0vj�x^;opX<=Av��� ��w�fwbRJ�����A��]a,���a��M�J�U�g6�@9=��51ib��0�w�}����K����if%c�c�p	�����j���'��������_���a@������_5�l��48�x���+����9�v�t$%&H �5�_$���|�� ��t�xi%���>/�ɥ�(z[�ԉ)�@	[��9��e��_Cy��ٽ���k �}/r)��˚?Nb̠��[�җ������݂�da�5��?$#<<LX!���-eT]�<��4�ʚz|��m�~з�y�9��^8�zd�λ��b�hQ!8�a��`��|/=�X�D�{%��]�ES1wj2SE����el#�V}'J���T3�6a�+d��X��c�E�/˛�*\�m%Ƽ�dG��J�|qEjE�r�d���dF�]�p��ε���PX9�����wV���X89��i������Hى��N�fqb�lFGW�j�e7塚��<�Ϯ<��c�u�J�@g���>���|7?����#!2hgC����R<�X]�(Px��0<���r���F\�I�:y8o�d����g���`���@�����[�NKV#9�E��`�-=�PJ��`j��A%v�:�r<�	� .�W<�8�M\���fŹ1>�Lא�����o�i��&��A��V��e��w�8�#tDE��0�[o���n�[j��x��Mf�iSR���-�NLJ���k��yǩ�>:� uTh �Z4���`Ɗ���<K�y��w�ԩ��D����~��a㲒��v��>3M|P�r�eu e�
�����H*q��Eh������]]������J5���Պ�+gG��Iy#=6 �fD�q?]�U	8F�ێ���]|%YV*&�����h����[���/?����K�&N�uw,�ؿ|IMs�|�����������j��AZM�[[v{fg���{7��o �H�_��,�T(��v����C�!\��\�s�s,a0�w��3x�3�Yj�(R~�C��/������"|H;[��7����gz�� 3;X�_��܇c#?i��~�����m�o����H+I�3�B�:m"�v����T+�7�"W��T�Y�(��}��A2��6#5bQ���+�g�صٝ�-mM��]��ܜ�����`���5��&���ge��>����-eM=A��4{�+�D���9{&��Ӷ�4J��:<^���N;~��YAnS�pzݬ��%>�ʀ�NE�t���*��m�C�V���xlN�W��f����֣�)�u=1##�a
A[�N�?q�&�+f�5��A�/��z=Qĸ�o~c���m�OuSN��F�w˺"˟c�U����������[�m�[�Z��
u��m}�0�@�b�k_Y��)5d8y�Փ�w�=/�s��~l�R��dl$��q7�G�����M��/�&D�vI�T���Q��؊�E��	
E��A�۫�X���w2�f��3m����h$P��� H�4��e�+K�.yF�sq�6�i���kv��q5���qa�e�;m�>zW����/3tJ����UM�Uc��s����+�A�fqZ ���tKcZ� 5 |���MF���P���__�%��q��ߎK�r��o��Ʒ�\e�[@�����lS��?�    IEND�B`�PK   �?X��) oj /   images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngĻg\S��=�2�
��>zSzG�w�BT���	�����N@z��	��^H'z �����|_�{�?~��疳�.k�}�1TS]��������\IQ���z"�k����Hg����\I�O��ߟo?���I�Е���������:�� ����������ks"OOOk[W��N�<�.��(	Z"���d��x�m�{������O��݇D]kg`%��1�hU�O\dq5�Zl��|�M��l?���c�0*M���Z�ZwN��a��j�ߕ��b���������ad�~���ޒL���~0,�Ƈ�/�7d�|��b)���_N�;��3H�xg���c�AA⿏eri:��>GB��},��i;�w���J����S��E��ٮ����G#�%�ܨ�1T�{���''=���']|޹U��]�b�E�џ?*�������W 
�_@�O㩤0͌����g��A)Z,��m��ąO�s��V��I�k9y&�+����u���58����|������U�J�t�ر�����M��/���;T�1yD2���k�K�%�$Uf�U3�W$��B����K��"T?ϗTa�:�
m�p<k$��W�����YeZ��<[
�7.�����5.����/���y�_���L�܃A����d+�̿��!s��!s
�W�B.�@�r;Ku�&bt�����4��E�Y)!S�!��,�c�����aAX�J����e��[5y���F�,����f�i��x�d!H��y7��<�_�Mv�N�Q椽�Ѹ^y��-9f�q�~�q$�W�
^5?�]�?C��5(��`I�VZ��4[7��|���H��[��S�M�_�ߞ�x"+P�
*w�M�n,5�p�?��}���y{�|y��omj��M�z���4ŉu[_��'u��}�f��!f=�J/��do���{�+��鄩A��bKw��|�1e�&V�~��I<G��t�1[ˉ)$���]w�ޝ�.Γ�Y�"pi�s���O��S���ſ�2�Ϳ6��]�F����n4JF�y0lM�C��!�ު�(�AX�o�֮�Ue3#y����ٓ��2<�`�;�C2�Q��J ����N��c�u^��a�&I�^7 BN��pJ�G��i���q��	�j�tǉ�z*�?v�_� 5�[���W/���)��6mwƌ��%-[���8�.��'7r���xћ!'6^�h �����g��NS��%gvu�sώ��.��7'$���J�L��}�S�/�}ٞf��|�kb�W�)��ء杜�>v�zQ{P�uoQ=�����d�ꃀ��b����uM���պ�X*���`g���s���㍋�G�G]��H +K��,�	��RC�T(��3;��Wτf1j��D�!�%4[l�w&�e+�:��zI�^5x�2y�A�9���7N��e����-i�w���[���P�Ն'lE��)$�ɏ���S��0�a�!m�� �`D1�װ(\o�xoz力�׋��D�߁ԫ]tg�g؜!��C���t6j٤��� ���Z�=_���c#�_Q3��}C ��$����mD�$~�-��I����8 ��Y��3( �s���6q�\�1m�Rc�B���Wu4~��Ū��h��2��z�(|+�q���9�h޷�+9[]�TS�vW��e�Jr@rB�g���/[a�W�1Z��������DeL���O�OyD��u�ԁ%2�(�����{�F��lk��L6M]��8�z��T�B3�x����Ⴑ���gs׉ߙ-�^�6/�r�O�CV�3Z)�]s�P�!:�۟����C��9j��Pa�2��l��j�b���Ml�	��'9E�v7>�o��V�1���u*!�h��ίޕ��	2_G����v����X����D^��l�I�YH����z�����Yr�I����g�}Ӫ�a ��c�Nb�wO�ݝ?j<������Ĵ�ZN�]`�
(��3�i%_�F�s�� H�U\�fz��kw6��w���fË��9}��X�Rx��e�y�d'-�� ��!��;��JL}+�����S�{9<���a�0%��i��U%/�X%��T#��'���䡚��3V�[��)\f�3�H�y�Y<�c��j%��o���vR��F�4�=��K����,�ұ��؃��`�Dim�i��b��nNT�d|@yLV&T�-<��|�K�1��#�����;�W�s�^���]p�髀K�ـO��.���?��� C����kLLH�#N�g��oE��NF���|�e�����!����	�W1E�!G�%�^=;Z�f-2f
�36��.{6N�}�S�;��V�#�A��އ�E7Hx�"t�t�m?<_՟�?��D2AkMb����P�Odv�.r���c�"�x/��|m��A���f�8qr*�����b�u�����W3%^L��[8�Y!Z³kG�7k~ز
�:�S�)
�����l�c\A}�����L�׵�o�Ε��`,���|/��K�G]צ��h�����g���s�f,��4��e2r��Z~�>�Do��6�C|v�g�u뛳��tb�CeOw��]�c���/i�t�L�N��{�7+?�pя�Y�o �W�g���u����&
F�fLd��o^����>�_>�����Ċ�/��Y9dg41���w���:J�B�s��XG��+`�<�vp� �Ê��2�&����!,��nw�P���ك�-�|���n3�{�����w��|:�n�Ȟ��i�~ʑ���;�l�}6)R۹=z��EH4�_��W��'�5���.��A컬�l��_�p�}�����'����ض�Lz�VΥ�/����ƌ���+��J`�hZN¥'ŐS�f�M�ӱMz]Ig�Y�8f��]9M�Ư`�SR�`l���pA����\����u���M��#g�!H���Sy��fm������CO�-�����y��U�&��+@e�Ǐ"R�1�4��T{{����LZ��Z�ж/��}���#U���m����:՞��g��ɫT��k&N�詝O�#z��"{!�زw2�n�r��<8�c�]jǼU6�r��r�>�J@n�W*�U,��|�i	a����˼��oB��~|I�X6�h*k:���݆�Q�G�M��P4d�3s[p�Uk���qc���X��ں���cCs�J�x�-R��tojg:wt��f|�9=�c�a��s��J~�RWs���E{"U�G�����t��tj�*��
��1ũ)��1M���ԫ.=��T�㙫�
����q���H�-u�H�0=¹@ؿW�Y1��JK�:�"��J�\=LJ*',=�g�G_{���I�~l�b��w��G�\��Vk��=�juڡq~�˪��:w�q.��&*XUz�"�Ķ����ι~}kI
�w�2�^��>5u��?5}��%N�*�@R��}1x ���4C+�c�����i�Խ��*/��3����O/܆�7�[_��W�).~b���������72�}_0������-Zluq(���*�Cb(!���G��.8[�~��ɑ'�y�#�N)Sh0��wЦ>��� 9�` 4%�	�m8+������� ��W(��Mlg��f�z��D*�-�ӗ������>t�5t�IO�]�v_w��DA74K��u���^m�1��q�6��xp�'q=%����AP^ݘ�ݸ�nt�t���t7e�Y����^r�]n�b�f��[�¡9�o
����8^հć#n�w4��*�}n(���r���Q��U���i�����8}k㟜o�ש�>y��,�;Ѧ��b�y��]z)�����Zo��n[g4�zٚ��ܖ��i.��[8��L��1�r
&p��{��2���/���k��G�I��%0R�ۘ]� f
�}jY����9�a%�2��]�0�Q�������k|�L��&�Txlʹ>��t�&[Y�ar�}˰�����F��q���L&������;���/WdГ��Z&��N��|�d(j��-b�r�^Cֳ����ܖq��V���|҉u�:>Hf*��e��벤�YZ�3BS�����|JQ��!�6;^G�#�g	>�v����L��yºL_�,N&"�����u�Q����V@�w! �������m�*1�S*,N1�g36�B��J�=2�o����/�
��L��}H�����\��+���������"NwC���-@*�+a���&�({� �����x\!���ԖJfc�ݧ"lL�J�R4ob�.��}���I�d���d{�DB\�l[A.�k�@����0� u�D�	��y�	��	w��[��^'�r���	�ƎިC���Y��B������/���P|��t��y�d��Y���)^6�{�:v@��t$��|�-�&.r��>� �L�zGjv}�	���OgFq��?6jF���)�
��::ߝ�^*���Fz��nOn^�8��W.ǭԂ��0L�:Q�7�<�~���7���t���эh�I��?�@E�?�o���v(:�����5���󼳈UW��P��Ʃ�8��~��h��YN�r�Mi��BNW\D�m}�θ��a�c���������}�)z�l�j���-��1S�;ǣ���л-�`"���$�.�x)xi׵!�rf�:ޗ�vhVLdc2# ������qiݵn��C����7"s�#�Y������lR�+�0)�Cݷj�yK��I���TgҮ�䮇'�a�׭=Z��ўL;⸕*�����@�ƛ�~���-�-&JL�ĺ1�bC�D�r�0�%��~�g\�3���=0�o���=}JEE�ǃ�3����'�/�p""mO�6K��((;;���ar�瓼�B�r���^k�����7���?�\&FIg	|�958*��Jζ̩�GV��!��8�v7�i�P��jɯ��z��p��7}/E�A�W�y����ѭ��D8e�S���1�]t�|v��w�v.`/�Un��;�U�P����2�d�����;tH\R�4l-=l��dZ��(��{��^�-��2��(���0��0��CF���������J�--���޷�_h�M��I�ޭ���y\ ��p�*a�;z�K�G���?S�B@&r��RC˟���v�Z�$�\v^��I�܈n�;[��W'n�~�@7�> �b��4�Kdq��[�2|t����蹃^��6�JRp��@XES#���?G��:�{�*/le�W����yI�u�	�~���VXכ��
����~Үk���['���1_3kO(h��4�Wۍ�$�ac�|�>e�  Ks�����'�c�6w$_p�1���c(�����~Y�u~��i)lG��k��&w��',���B#�ё������m�u��D�!)�]� �>�Z�2�>�fM��-���d+���v�����+��(��S6�X�B����"zLycC�рLm����7�U��0_��l���~hH3��N��JD��1aP���}[z�W�^x�Rt�;��<g��2kS�V�g���W�yꞶ4v�;�\'��w?e�۱�]C��{S���17�Q�L�����	�Ļ�y��\I�y7F�)�uk����X�D7׀K��
�yQ
��ρ��rXpm[[����$|<{�ߟ��:�S- ������� Pe�'|�uF�*:�"�6��h��6��w����:��=1m�ß����-��"7AՕ���Q��/��s���ve+�/JԣM`|��f'��@����� -��͎̀����!�w���'�$�>@:= ����F�Syy�3��D�\	���C�ʒ3�� ?_�U#���g]�L�2��n�~+}��ח8_�o��a*�X5nSD�w��s���g�"��~�i��ްO�mLs���l��}�WyV=�^���(�*��c�Yy� g��'l�Cl�M��X>�U�.�\C��+B���hi	��v����{:&&�[ȭ8UsC�@�L)�P�6VV�<��Bm��y��JߑXXі�`x^Ͳ�Ӑ�~���x5Ke�޳;�F�	"��k�BGJ�,�\� ]���b.�aC�ً.��s�0��r{_��8[� P\ķ���������ʠ��+���f��k�a�ݦ��!Q�⏐
�pAMދr��k�&��%3J�7~�%��f�n���ښ��.HI�U�@`3�[���޷~���9Z������{=��۾�i�9�s����k=<�7���8����;�!�~����\g �D�筕����~^ѧ��{��"�H)l��h��O4~|�n��?��d��a��HU]�A���L�k[�]���_g5&�V�q_�|��S>g뭿��a����U�����9
���vp={��O7���u�ѯrarّ��ѓ��2[%Zmk��_O�l6-2YTD�f�W����g�+�q�w5�~8���8�nD]�V�Gv�3"9�,�M1ar}��m��E����"�{Y���Q����6�U��U�,ܒ�#���t\�dU7�`f��ҫŴ����0Om�e�:77��OC����$W��=����x��{ �X[~�2�f%�8xO�X�[��-ADV9o��D��%#�G�\�3�LR\V�c�N��}������Ís�RuY�\;2Tb�ǚ)��3��V���I��
Q��'���5���F�&
��$'8�f���A��ɄD�ۑs�I'��𻛺ƵVJ�M�?��U��Ǜ'�1Hp�<�Rݠ�U=b_d���)�Rf_�L%|�`�=�]���,�+��G��&��F;5�,�Z�I_X+q�Ln��ޙ�~�|����vT�5�S���v:�P@皂�V�>ݞI,Iٔ�"��%塡ɬXNgh5�w:]ۢ��A��*�*����Z@����H�L�;Jt� ;[ ��4m���N��6y�U���kq���7��������8��3�m?l��'ޞ���j4���g���b��s�U���97�|���`�{���2�1��]L���)�6��k,��Ї�:å�ۂ�<U\*�55F@�3Y�_\T�g DD�a���ɋ�����\^N�.	���^0�^�R�����L�c��9��S��I��}R��ӭ����iX+���~�n��˵�
�/c5pgS�r���9���e2��!�=�#��W��j������r�]|��>Y7�\V����ɪ����[��m�J����u� �r��@�1�6�1�ĦX�<��`�e,2!~d���ex�b��`�ܨu.�{�h	�2�9NN?�'�S^B���wGa���3�9��ɺ��PBo�9�ae�Z�^8�(�``��e� m央�Q�G�T�a��� ܌���Gg]0���^!���k�+�U>�kvWx���l)��&�X>��j��7��e&�<aw L������>��!���S��B�m��G��>!]��ʟ�j�o/�PQxQC
e�/`jS	?;l,07P�5��a�ѽ4���o��#P��bwȂ?[�l�q7P��'H��G@���_nشS�FR�ZJ�[v�vO��q:@��u4��8�3�4�z�f�����\[S��\YCW���0T4z�-�U��J.G�m`
m<����e~LoN4 1�����5��j�pj��#j��x9w�C#SA�����
K-�xN�.�K�i4�o��(��D��٣���K �dP��Ј��{6��@���lʞË�7K��*����@������'������:�*�mp��^���L���Td���
�u� �n{�f�j��)�;�d�4��Ƚ��6MQ4�
AO �|��\ݸ����lD��ig���o���Tk�&�S�q�ǌa_�p��Õ�\����d��aR$�buچ��]q	,ݏ��4�6�5އ555��&`�@��8>�.� ��>�N鮸i���Y2�iP����c��<���p�l��;��&Ӗ��=�	�EB�C+no��Y�ۓ�<����J���*�l��_P�P$j2&Vr62C�ѱ�m�Ĵ�d�ׯmn�~��Ͼd�Y��I�w���H����ۃ�z	ey
�xYH�5AIM�<\�J�Bi�9����SO2���J���u(���U�fC����4�]V�o��������J\xL��j���o��wg���G���tL%A�X
 ��f�-�]E%wa��lq��9�ҿ[���c�]�� 8���I(5��b}c�4����/;8덧�G�џj �~+�6��?�ߜ�,]8�Ձ������U�MTd��;F �$v/?��&t�z\�2@`q�|�?�g�.����Ϸ�Y���j&�%����yԣ�j����F�Zw��C�������c�-[
+�B�aUE�S�<~j!m¦�Wb���j�уy�K�vΎQB�_2���H�`�|mh�:�^���zA�Զ���f��Q4������|���<Wj�o#���zNm&��	ͭۻ�k�����o�x�=��N�pz:9�9Jh5�=����&H��z\�����X��1��������s�S�rkF�	K4?��c����]ߜ��˝��v\���ޙ7s�\���#
I��SSu/�7V37�f��ǣ	���	�U,|'Y��8kd?W����������+ ��6"�]o:<�]�6E���+류�I�q@h���Y���{(U-�ʤ�ؗ�.��R�C��q�s�e���"�xr��/�<X��.VΞ�6�����|����%�\
Ҿ	� ��O�����Te�X��9��%��x��녔n�i[�)���El��4�����[��u��ae
�SVSX9��<�Ǉ��,��	{n48$��K�T�G.�D{{�k�����k�mG;��F��|��2i�m��r!��N��2����.��?-�a�C�s�,�d9��y���G�r��6ڼ�>:w�:�	`��H�Y����l��#��zxdZn�Ď�y��X�:/��&���%��0��<X����RW����s�yK���L[Q��/�ϛ4�6�-_�4W��蓡B�>�ΰ��۬��O�QI7v��fKh$�be�����ٺp��z�����WA�)�����vH�h'������2�bz8�F�Y\
���wv�j+ʗ��LM��K�<d��l	�j��ى��C���&�W52�"�J"B�'�*-(��tR�����р�L���5�"�~�'UjZ��j1|9o��dT�T� F���P��`���.��e^O��Lk���w^;�>�*�=�b�����+Qn�N����Z����&#_��oV/��۩���νKZWrB�A ���w�b��I8{=I2�Bh�MM+��vu���8A�ˉ{�δƓ��!I��풴| e��U�{��Z�£+��@��o��B< ���H���K�s+��R/pn�@�-��cִ��\W:�W�x����=��e�1�g��Y1~���e�$'=~����L|�d�|�~�/����/��̘V[�kmCKe���r}s��_ӥi���+�م�Z2H����v�ϒf���g���b�V��0���H���ݠ�H`R�`9���ۏM�o�z���,U��%G\Jt[�:�Ӧѣ�e5�0�{�Oj����7OJw�u��8}D�X��(?�d&���{���`.ğ>�;��Q}�f3ͣ���&.)��#����+5.�J�A=�o��o&��,V���Uߘ��5*5i�`%��v��z�;Y���C�Nf�D��{�SV9w.u�������ĝ�����f>B���^��c�����!�n���O�*��%8�UO�������S�'��6H�,uO��rG��.]�t*����a�_8����ky��j�琎�
��7�\���/����_*� �o\ҥϊ�s���xr���!U���0��������,�`�.(���A8��H��B��*<����]2v���f�R���t����*�
wqO�F\H_��I��R�;W&�g�	Cq�,|���U&�f�=�"�݁��W13(�����=����!*�z�h�I����Cac�Ϋ�m�C��3	�Y{��@]���u���������LWZ���p��Yc��;��|@l����*�/�*VC�v��[��)Z�`�ӝ]��y���׏�ofl��e5��d)����PJ2���󰜙0���Y�Mݳ0��YQ���㟀�^b���|j888X�ZJ��&s���x�P��b!f&w��a�`��	v���}��](�q��<Sx��t�-��
��*�QU˲�]��ˊ����W@��dq�]ۇ�������N��T��ap����4a{$#��ʵ��#�XP�<$���#\@�8�-o=eT
���Ĳ�C��FNx+�+֓}�)&�M��/���8�ш+�X�����!$j�=��{�G^�_ NN�~{5���R| Zvg��	��Q�3�h.X=Lf���ߌ����lQ�=��O��ٚ�/o=���ӳY��,	�g���s���3�M;S3�*�9bS�i�>�OH����3S�Q��R%�vdw�1PX�.����oD�D���a�,�g��l��U��IF����5 ��}N�!�R�V��Չ%��c�$Se���Xy��i�}B颋m.��� d�2U�m���#�)s%�}���ˏ�O=�u~�z����=�81�$�1F�P̳267�3Se��1�,����0��'����䖅����D|�(�l�?�f6�1�����>(p�.����1E$G�<A���p$���t�����w���QNr�nAY��s�I�Q�)A���������F��i��q�H�\+�wi%9n�'qU��%_:�d鍋;W�c�?�q�5Y����k���c	۷����t5ޜ�s ����H��bH���Ÿ�.���Ƈ2�x=��zV$!�{C�r�y�� \��<��{c�_dT���	°�ժ;�py��顺��.)��םO��b̊�V�Yn�Z��0Wre#b$N�k6-�+3��?��%�*��d�!8UH]�w���z�ґ�Q�L�a��$�T�A}����E�\ �Xx����?C؁����bM@:�}����͚<�/����`d,W��(��^:�s�	i�V7�1e�\�c�l��G�
�˰𓾰&��{Ҁ�q����^�48}:���j�=���X���3�ڴ޳����:l[���w�o-]�����i�-T7f�{�t��~�M@g�L���ä������+���(�u�fվ��2[^օ���{d�Y"�0����I����!(��P���|�IҠ	���R���o�~�Q��,�4~a�c5
R$�;�{������Mռ�u�����Z5G�xE�������a�/�?W�UIy�#����@]Vb�����B�OK� �/�����6�ɺ��<x�d�@ �Q��k
�Nv.��6�Ȇ�r��t�۽؆��u�*6�YU�_fk��������C����Q+����6�ɾH��6=��Ǿ���'3rvWk��x��O�.���{,��{�G%��C{.���VF����{� :��_ʨ�J�#oPo0���[��HY\��i|(d��+��8��D'�PKk�Gٍ�jl0����2�ڱ���a�C��Z�km���&�}Z�?��v2�>���߼
~��5��g�;�#P��M	+�1���9��z$?"����΃�M��/��4�{�*.�Ѐ�����>�S���W��I�wy�r���y�^�M�K2 �NP�q��!�Th��͟X);��ʗ�H�`�<ᐾ�[�i��'f^�#�R}z�(���/kE��)7��$��ׅ<��[)�
�֍CJ֖��'��5�3�j�lPs��K��V��aO���l��YO�|��O|r�5Ua; �H�-z�a&�W�sH1�	+�#&~A)�m+�vD�%�U}��z�mN�u)�z}�l��
K=o��_�_�?�OX|��ǋ�`��ir��$�c�]���_����k#��h'���	�eS�e���nB���4�&#1Vۍ˶��I��p��ں4GIC�kc���C��c��8'��b���`k���������F���.!��N�vM�r��v�\>�Ą�7��M���w�Y�f��v}��Sb�'V���͒xp�!�2xUU����a�~V����gxX�.5�S�?����r�5~)��֪%�]{�+鼘�7Ӽ?�Z����G)iTOb������������(.Y��ŋ���P��dڬ�n��{-�	cݜ3��Z��3�:r��S��G��2#W��
��jk9nF�Qc9��lR�]�����[{Ψ�z�?���]4|p2��`EMbI5�B�+7u��fɝWР&'iֳ�7���bl�����<L�E\#h^=��B�����_��;���^Y�)`��6d����֕^����r-*�j�)��p����ϔfH}=uH-����2Ϲ�$&�Y�x}��\j�F�c?ơw�qP��nq��/���P�fs]��.����ݞ�q῁Qӿ�;'�&t���o��y���6���|��X�p�1C�އ�K���9mK�����P=���}_/�� �u(�8/ƼmNV���t�D��d�ed2M�k�0���O�N�)�ք� �ɫ�k���Q���M���js	�vU��7��b��4Ԟ���#
�Gt�B]��o�0OOx���M{_�3tw_��w�`�>v��/w�it���J�N?�2���	�Zi|�:FR�����7`Z`��?���*�Zn��F��~a����{8�X����=]��#zh>�����Ԋ���b�Yj�#�����g
.�RQkB?.����|���]p�g<�����֓�׬_	T������2b!C�E���x	�^�U��/���m�j22gՕE�����]�B?�B%��J�$�j�����,�`���}�4����<ӎ�Z���&O�k*TՈI�] ��Ӟֵ�/XA�=�[�`VN��f�"<���S���ه��b�w��`2��.�X�7�Rm�V͑�Qn����V��x�G�������o����z���|��I�?�(�ܙ��¯t��OΟ/h�ǻmZ�.���j���?���*�%�ʟ�4L�.#���RVE�s)77Y�s9����? �io���X��%�-���x;q�p�ˣA�ҋ��v)?
)᧻����Z6V0��\��;k�( �x* ;NvT��_?=��^3�xЋ�*
 (��(��m0��V�1���)�G�;�Տ<���t��'�m�����a]�|�hq^�N�	8%���Q��Ur�SF�=J1�p���H�0��m���o[5sg[�0������_���^�뽿�_RV��u��	?D��U\���_i���N�0�v3�o� ��~�ɼ�
AR�;�]�n��?���
S�N�\�
�vt.P���+K��?�_�xnb��,ȹ���b�;y��f�����Uǀ7��.���(����HQ����ôh#>b��u]L��a�/��fx��"��L��<��i�!N�e���X��2>� ��V:��3v��QB<���������A��z����!!o�X�\��_hPIE��Ѐ0��}��Gf^}��%��~�W}D�v��t����#vy�Rh�?_e�*�Uv�8Πƞⵝ&1S�6��D���n�$��F2�׳�Gقz:q9��k�3�:�}9Φ��>fmL�M@�V8̏_*U���?�;�nK^��y�-֤�-�:	h>,�w�K�Z ���}iwǡ4Q
u�K���%�"j&��t��O
�6�����v=�8���]\S�HŔ��[xzڂ��[ג�H�$?�Hz+��$����÷�}yt���WC����ؾf�^E�+��Ÿ�j��d���i�]�I/j:>�H�����3�B�a?���ۇ/z�k�:M����N}'���6�<�M{�H���x���.;B/�r"��l������O�c�/�H5OqzJ;�|�bSN��#��0ʺ����z}3�6Y��y���\��:�L�Ld�O__j\W����"WWwwrt�"��3�B�����_V���bV�Rb�Ѽ����)����az,[]`���s�}��$>~E�R�=��=3�޴���/~V��e�g�F>��]��'�MM���Y�|����^ѧ�Yeoʸ:iA}l�OO���~�uB�9_�ڊ
�r����I����ݐ�<��'�w�n��?���=�}�U���EH�%^�D�4-L��NS�%�Dg�T~��6���b��rl�ê1]����R�5/G�#�O���B��vy/��K���ϓ�|+���S65m�!�37�S���S�,�3z�
4p�Q�]��!�o���1��-n�IW)�g��'�|���'������{<��W�U'���K�1���k���kc By���� ���KW��ge[ճW����=�WQ�e�M����Ǽ'�Q��S�����mUe���@�+��ѭл俆�㲲�߸qC�g�q�h��o�ݏ�%��Q}.�T{�
�6�R��|�yk#1#����c�W����.f���Qr~�����}w;�n��\$���=�*��`�2���C�-��x�:)OjiTd�"�>,�}�_H�����p��|�������~V8o�6�^�u��ߵ9�~�
m�=�Xn�Pm��q2xp��h�霺�t�-��}_�}<;"�W��$�bl�q��-�E�dcs�rb`\�󮔺����8���^B�f�.�Ul�,�>�����{���\�ԛ���U�%=Î�`w�zGH��=����8\�2�?cgz�Nã�tx���_i(��ݩ��g�S�� �τ�+�;���P�	n]�ҧ_��6N�9a)!�mu���k��{ɾQK���ڗȑ��DP���#��I�^��b���T�{�Q��[ʥΟK�d��	�h�?���5T{,L	�N�GG~�brS�\��w�xyҼ�_�����F�u��4~�	W�A>�����R)�_ZM|Y���x��D��4��C���N�>�S�ӛ���.���wo'�<[��|֥]��ǁ���<M=�[)�ܙ��.4`L|�N���U��-�Z�Bҹ:{�TGa|�e��������vά�])�:]r�p��3.3�3u=>� ��{_,0����&fͻ˞��&%�/�����!��������D��o��a���)���q���j4����	���l�u�$fZ�_�+���eRW�|�������0�����sc	��Gb&g�q��3�t�򛿼�Wi�7�E�b��$��;���r�U�b��{�*Skrپ\�m��i�u�.'>�0�b	����',>�0�E6�|W���6�P��#�[�%4�O����yX�����2>k�D�<�����uўs�
?�.��-�����t>x�h��rҴ��a�f�)HY�o���;�
ϑx"U�^Ys�H�;�-����C�<Ðk�B\VKF�Ya�]j�u��t+��H1|��i�<v$�]4��S��U�P�9WH�?sn������5�_����bO��~�n�r��jF?�_p�`ۈ0i,w���`[%�����������r�vڤ��y7F.�Ky�N?��c;�^��D����<�� �k�t��}gZ|
���vv�8����߅"���N�_�^��b4j.42��c7h��CL5��K;�ɣ8�w?�u;btK}*��O)\цBu�c��cz�o*N\�ku�������3��F4�?)���ԇM�f�D��O润��')>ʴ�x{5���뫍W�4��nL?�tq��#�6�i�xy���49�}pP��^�+f?]#u\���s��a�1R��'����x�~ay",�e��g̶�'���;[�S��{Mo�ɀ�df'���C�\ӆ}J7�����Ơ){��[߲l)4�s��'��)��UA��ύ@��JAb
����b�
2�ѓ����q�:oi^��y%���q�V���3�Xv�n�^��_��-�1�!���͸��^�P���e��V����n)(�r��w�k]|t�mdP��>/X74B[;ܾ���	@� z�z.Df�}݁Q���n��IA�Lg;�����0܀�9�w�W�X��%#jv������C�aS\�f�������hi(ɯ�Q�5��6$)4�|~��su}r����Z���<r������י-g��F��_B;v20�ߚlK��E
>.�wS��?}�,� :0Z�}4�� �\��)>�o������q�㤥U���<�fX��¨�K��[r��S꘥�ƶ+-��1:�s}����h�(>����1��P'��wa�s�����q-�JӍ��uy�t8���$HX��x�P�o�7�k�U*��t)5�o=�#���Uǘ{������^dOB`n�����3\�� �ڶ�uZ�v������9���c���w��Mn�
�J͸����]܆
��^��7��L���]�f���n���C�[��
���!K�����C�y�|]|�������ѩ�z�5�.�ů5]̆w�)��[�xa��&i�[=����vW��[�ǔ)�{�LX�������\��M{�_�=�sx����F����5��!��]�ݤ�>S~�K^��u3r69��5ɫ6�E=����mv�[r��V+#1_#7�����J�1�,�UFD�ȳ8�ͨgs���=&&�}|�9�w;�Ь�ƽ�A��hR�K-�n���E����,���Em��e͘O�>P����{�Ze��?���q�<���(���f�q0�KV��Q2�����]1'3��K24������$�*6�c"V��\�SέkG�-wwhQӒ�����xX4�,��V���Ӎ��Am^��D���_yVj����}��O[,��1%�@q��Ɩ�Aa��Q_�����y�;~�_,
/�(8�|@`7L��PW��@��;&w��^t#���,��<(��h(G?4y
�7����Lb�I��S�7��(�_+Z���F�0\�ch���z�xc�=���k�$���k�����&�A�CB���A������S	��;�����Y�ߢ���;���0�����\׉*�ݒ��ް⛹6gv���5D�bO�!OҜB�߯�ԐT�B�\߽�l�ȢW�[�Q8���Zk].�p� ���\"�G|Q>~��s���C���Ć.�tD��;����.t����\|������d%N2��4����WxG��]�7B�_���4~���ax���!��BZF�}U#����wϊ7ڊ��s��wM��[NԵ(ԤiT_��4�$���Cr;����b�W�������B���?m�/�{��'Pܕ6��~e�H��{�۟_��L�Gpۂ�Z[��z�YD µz�hT㲷]���b�v�Ma�T�M�9���C��C�@��c��J�KY��yH��x��-�h�\����˒��m�8�r&����~�ގ�j�G�*�d�qB��'^޺�M�X�y�f�Jg���-y�l��5��_���UxU��9M<�	�f��c�4���I�V�!V����`��"�B>ka�-������%LȬ�h�S`b51ӥ�y�7;�FZ\�
�#.�S��Q2�� Y�k�>���@�E�����__���}.���Z��{+�:��
!W���͙�(�r�Z�0�^J�����/\[P��h�lR?M�
ZB䑬9��8Y�ۚ��w}��E>�3����x�8�81��wQnn�i䷱u�����z޵�3�Bp�Z\��e�RP�0�tw���8�y�t���K����7 G����x����)�p��B�q� g�;������������Rg��7�w*�]��!���?��E	_��t���j|R���	��q^�6o��SΘm�5��r�(<M`�o�s�r�!�9&6��N����+�{Ƃ��K��N��Y��5�CfL��Θ�G������b��&��]������qO6��GƧ����e���U�ϕX\��>R���p�NW$M��T������>���ړ��L��@؅�d$���Δ�Ҥ:W\Y�4��m�v�|`�[�l�is��)��*�^�����+x���%<%g��{����D	v����Y��5!���Vk|>��c�?�q�J�I�q쩕�㶉%���������^�*a5h֨}u��)k�yc����0kv������ <�$-8�~��پ�9ލ@or�8�fCH*�l�]������`���1+L�xk��M��u�o����.����?���8��w��m��*.�k��	��[*�*R�������v���bv�Lm\�v�	��熥����wϖ�ֽ�gZ-�M&x��*�̹�9m�e�.Q��$��l4�Up<v�f�4ġ�"_F���-�)v֑2�C���/,��0�������zRy�ɩh�6'\5�U�V����IV��!��@�����l����Y$+��`�ݪ���{�(M��Ϙw�wk��ri
��~��K�����\���T�����v�cf����e`��D�\�5�I��z�������8�{�co,E]�<��o����S�X��]_%�_���$����D��f���̂�L�` ��?��з�����S\�d��n���ߛ� Y����*6h@/�{m�-!J��~�
5l����g�m��ւ�c�7��[|&���ה�isC^I���f���}�#�hHVr�1w��zgf�(Y����5uUf����K���q�K����u7n"�V��}y�y�}!�'��������4��p-wخq7ܬ�S��&އ]�UP�~
I���x�jC3�z'��y"9&�Lb��e�V]�]�

���$(l]Pm�ē*t����sw�ur���(+W���M��*|.KMQL�@H�ztw7R��j���mӹ��Uƹ+�K�|t
@��t ;��,'� �n��2ŬKZ�kL�=��th�L��\嶕tt������%[�������VnR,�'�q�)�̟���u(���b�/�����sr�U_K�(��~3*1�z�v��l��c�s����o�|6)�~a<�Z�F¤������0����Q��3����鷙ߪ�1�(���A~��B>�"�~2�[.onU���;~\ƭ���u�Ga��l)d8��ψ�I�Pۖt���\�3;����r���vb8m�7*����Bzi�>�4�Ĺ	�65����hZ�AZ�ڑ�#����ר��n�KJQ���/ú�1O�'F���!������ �781,��.y���F��:S�"(����8>�����''��-��3��Jv"	�k�ר�֗6�.Y�7�>/E�N�Cg�&��9)M�h����L��[e5���q����?�F! �<�g��c⡸c;>Nd|�:R��x��"�+Y
�	kƬ!�����k��n�޵����-�?�;�@�ԭ��k3�x�ѻ>��u����b"Ԩ?��q�3H:rݷ�upq��È�����x���u�`{��`���q�:���he��+�Ն�,u��c5�,��US*�Ō�=�r�0��L���љ�N�֮��/�o�"����� ^f�]�q�-f�tl���5�� CM��M�NET�Q��T|#c���@FN�|4�O7��QDDDp��gL���=��gޛ�I�ȵ"7a������%aI��2��O6���gغ����a;�U�9���Q̏If̋��|���n#�}�Fϰ�%W]��m,U\���׿�������mV@O[��é���g�����D��D�wEBӿ�/�`��A�G������K8PgS�(�}��)��..�Ws�^������[��s*��q.[�����	����ݮ�b�cB��Ҋ	�>6����]ە$���N�[�Ǽqm4�#0�S��Y�ed�44�rhY���*�"2;���	�Ф������Cea�}�aRO��a�0�F��:X?�s��R�?i^�9�����@
,{$�z������S��rDiހ(�D���50w����N%�hE2@g��2Эwa�!�n�wΟ/	eu�ܹ��_��O�+�cBvU���/��1ש�_�;�� ��<d���/����g�V���Xr���&���У�������M	�6D���.��ll0��C{�?竭b҅���G��-7:�4�?u����S�ɷ����HQ� ʄx�|Z&u$EY�TN}ϰ�CRB��]̬�ٵ|�&lw�vK�S�6�k�zʁ�r��1vG��eҘ!T��ӑ�ɞ3����Q=��!B�nZ��vZ~bL�ro�q�v]]]$����3���M^%��{X��v�������)���k���}/��z�G�Z�4fu�p���72�]��/ ��'�Xu#3�P�)/q7�6�"k*E5��/p���Gb���9�y'~IE}���:X���ڨ����;��X�W��f�p�ՙ{~rZIӷU�j��)�J51�;mo\o��R2�Y�{�xR�V�����d�YWiQ��vZ���F�]頃�UB)��ue�m���!ϚC!X9Z��3c�y�?;�r��;4���o�gN��ܔ2�T��?63���-uBu�����*��mG�����r���
��e6��)ϑٴ����ǂ�F����|���]8��%`K�%��ђ[�O�V���^'���8���w �J��Ȧ��3*��@�S������RD���� �˒6+u�����T@�%2�YC4\M��񢢖IJ��C��\��e5a��,q��]�{f������&=�����*\�/�1y������Nx�sVjZ�:2a"����A��ba���|����� � ��UQYp����r�������S���[�.2b1��;e�M��{q��z=ߟ�a�l��*��^^���׶Kx9Ԉ���W����$�������������KҶ���M+�����.��p:�&\o��e�?�����|1�?���A�|��(�ZP[��P#hځ�c_���ٌ���ռ��a+���ֲ�?��!<ɋU����D����Ђ��p˛����kt�a�ㆵʤ��R�,��H�	��Z��8����g)�)���JOx�P���n1��ف&�$)Vof6��+�A܎�?��|�P�2���ԋ+�n�Kˊ�^��/�_�j�}�S!'P!�Xϟp)�tw�Q��Cx�S�d�j$��i���㝺�h��N��� �Y������ۏ�m,�a.=��N<�XЌ0�54�}����{�L6�І�Q�^_M�\Z׿$|��;}��N�0C��,^͋�k�C zgW���5�)�j���fl-$Z3y�(tFT��k���!�h�2&{�9-2�����1'C�CE��u�|��gE��x2	"�J)���u��Ξ��;C�Y��{'|l={�,�������%7�Q�c#˽F�9cw���kɅR��/��!Rsoǹ�/�&ٳ��!\��X�#��f,z�s���/�Y���6�5u/:�[4�,�����E��-�.��d��e�J[�ߓ��܂^b��O������:y:���O�OgU�#���f���4��"�݂�|�|�7Vi���w.`6!߫�rl�m��賬�{�bI��"sB�y�hȆ$�?�����"(�޼TBA]`�X��/���,b�	=�:iq5���c��hږ I���y^� ��)�}�^���?���L^��zv0�z�DN�<{9vv��Y���u�aP�ƀ���tdѝ�1��ތ5�(\��?�h�C3g�sM�$��C?a���
��|��hG����{߿
���������w�w�fo7�<�U��d=~�r�V6�i�� �V�c�j�^#�#�C�
�ʑeJ2�r&����n���1�'`��z,]��A�a���5ݜs^U-|_�G��b�p��y)��l�4�&�B2�iQ����9}!pS���O��=�Q���Xn�D��,��o�z�[�]TRs>����z��/U�����+ދ�>�������ן�8�ޙIƸPK,�3P�#�1�m�i��=?�H���"�lXC�O��R�x��8�����v�_���<���:<I-��2J��^e�(�O:a��;$8�:�p�:h�+��<o�C:f�,���:W��;a�t]I#���A��{C�/��й\mnY"��0w[: ?�s}�9�,����.J/	����%����ӵ0\��WN״��ǿ�^q�6;D��Y���/�9����>q�R�����y�UJl9[���R�B�L��X�~%o�Pgi�t���;{Є	�O%nud�ʲdn��6iC'�c/��n��g�&^}_������8�/&���(X�����2�H�Ȼ\�O)����y�1y�|���C"��eq�L�5S�������.�����?yx�Qq���h��d�Ui6p]N�mQd��o_1z����+�vYJ�0�u�[�i����6<)���G�2v���� ��`2O�ڃ���bÎW� �F�y��&�t��DP��c��Q~2�rDkb�͞^gy�Г4Ѝ�*���'�[�"�����G�����@=���܌��D��6uT�����z�v��W�>��_�$���IY�_�~�P���>`�u�p\����&�v����%ܶÇw .�|̃9�~�cBw��U6|�,�a��ئXWx�f���(��>݄�gOl�c�wO����ݮ�&QaEY�l�!��k��?[u+O�A����Vv���%C��Y���'���1AA���^$%{�W`���sR� 6���hpm���H�m:����j�-�j��?���dz�;�#��|�j��ZAp�!�FB���z��3�
�
ae��fUb�z9�b������S�cd!ۛ`���<�v��=��g�#�.�n�f[�OΙ7u�G�f�.��#x��=��������&�*�+ⴠa�opa�,Kp�E��m��ߴr<��8r r�SY�\��tn�����7��v�@���~�_�4�����֊<���3̒��WPN��'1c4
1��TҎP�Vf�]��o�'-;�gw�p�с��|��_�nY�}0~hRme����ѴHڢ�4� �ǭ0~{H��/�|1a�X/��(��T�I�s � �
1?�k=04i@����]~ƚ�n�,y۾/t�V�f6�.<��_a������-�z2��5���SI�Zx�z���L%�0Zx��%��F<���;��9���� ĩq��J=P:K�$�|V�b��z�6v}%�ni���X '�~Bp�.��'{��e.ᡝ��{|���e��e)3�x��SY����HWb�u^*��|mJ/��ǣ빅�53T��cc"�Y�RQ�!�0��t�!�-��<b�"�]0��_.�9��^�֯'��$c�^�u$��)l?�IN�5�?��.M�S-��ȣ7��Y�H(��9�01���M��:	�c�����%��Ҙ�h������a=� �[��߽l}%f�(kF�q��P�hq��f{. �M��d��"|- �/�k���-Ccq����(h���W�A����`(Pvu-B�a�k�Hxۻx 	_��+<2B��ٿХ���"G,������>��n�k�ׄ�*�ί�0���U�0�dwz�BH�?�-j#��rr���/�C���}�&{�㵡c;hB�	��tȣ���0a���\f�L�܎�Ƈf�A:�=;=3�������>�4�9�.fgl"�f�x��賛o�ۙ�F�~��-J��F�>�6	���T�����B�4n<$�_=+YF��\GxN�L����pUPЁ����p�����>~�8|�j�,L���~�^aS4YƆ�����'�֡�Dg��3�WHX�^����Y3�[n��1�"n#+�Z��׎��H�(��d�dYfb��2	��&��u���Ls�i��1)Vzd�2�s��d��/�>͸ل���r�0��z�������������F�9�5P�~ʟ%&��{р�{�Ӣ�˥}��~�4�u�8tI�U$����~�m+�-�� òh�/�<.1)���JT���L�P��|gRAv����m���"�m:x.l�B$b4:��t��x^�K�	q��]>�Z颎�/w�g����̩U)���Ƨ#�U�17R��Loj��/mz��YG�������\/�N.����ӻ۝����K������zOd������￉�%�M}�Q�p�O/�k�����A��u�6o�g����~T�a�N�VI�b��"�Od;�Ϯ� �w�A�G��d�����/��ߠ�F2IA{��V�2�n���jtzU�{8*�2������iK�%J}���{2�{g�#�@u܋�/�'���)s���d-����.����V�д�����ZM�9!<:P��t�>=�w'����A��P�� �D����R���d�k�
��31�ܸ7�"c�/�G��TbĬ*m^�R�}y^��LL��f�'K�И�94�P��"�\��j�O�_�>��a��tbJƄ� ��Ij7�t��@�ko;�pZ٢�6�*56$�����*�U5�|�O�o���5��m\���<��s�5��n�?2�Ni����EG��h}�|�����3�)A�/Q���Ң>���6 �l�tx�1$�}������c��IsL&H�A�"Hj��5�7&��o7J;.��;q���M�2ǧ��{�USB��'�O�)� �L�Љs�ۓ7�I�����d=�.�d�����5�c����ِc��c�7�8�Kē8�\}�����s�ګdA5`���8�c?���>�cxJ�s�6��e"�_�$��ޕ����Q�Z
8u��Z�'-��J�#z{%S*�0����M���ӕ�/�6�4wuf�툦s@)I��/�{�	�)�z2�S�j�^��d��\~��A: ��$ʺ��׹��tX���l ~�]��\�}F� �ǚt��6�;�V�xED��8%��g(�Y�Puul�S�������&8�ݜm�2�0�N�vm"�V,���r�L��u��]�Ѿ�&�\�ox�O���Vj_�|k����$	'E[�$���@<�E� ��8���H6ϕBl==���O ���I+[�LAG���s�=��;��R�	p�f\���_�k4a����bu����M��6}~M<Zo��T *L����ex���gT|<+&�v���-��(��0n���$����W��"%�'1~I��bB�ܑ��/Jb�N/h�ܭ��˿�uzˊ�uS�!0qh�i&f�"N��=��5H��K��6a��B��=����u�I�͐!��X8N�p�ȳy���!ȋ�Ȅ �
)44�&?�c���z����+�7��.�y�c�x�� ��j�����H���5vu�t��0\��\�5�_p�,4U�l�P��t
���(Y�1��{��C�S�Ab�G��5{���͑�1�r���$�'Lں$�b��s�v�a���H{y��/7R3�k���ٸ���>R,a�M�8#un�D�Ӳ)ta�-, 9�:0�����U\ܧ�:��C%���M?�$M\?i����u�˛�{wD܇-���C����giX������v�Mޑ�GC�����2%�W��m�G��XnaGiޚI&�b��2^vE&�P�r�dn�A��":�u�gJ�f���q	���q��.~��fQ���ĲTZ�r��e.Ј�LB�e��Tv�C���7��ں0���|=��s���.�.$E��T��z��vӕ~�����q�=��A��v1E��[�g��\�&�̐6	F�_���Y�Bs4{/"|�x+5��R��*�!B�4�Q��l1aP�s�>@<�����^S�gS˔�TH�cD,�'�ٙ��^��ۿ�r/;�?v%	�a��Ļ��t_�z�^�E�%����+��\��'�
1�JN�R�����Ј���o���yqWG�&� �ԥL��)7[�g���P9�k���'�ع]��6R��H؀:\VD��s�` �[D+�+ށxc_:.^�jAPƅ��$��*h܁,{� Us�W�u�-�V�~�!q����G�N��{�9	h���u�ϕW*��YHrH�m�PU�I2�}���^6��m�9��T/!����o��=�0���bb7C�����j�� u��lO�3\!��M� O3uu\g����d _��O�P
��40���&���9B�P ��w����㦃���R�|{�^Ts�qb�CF�B%z�_h��1R6�O������OH��3g���1]WPx�n�JLsH����Bs��[��/~��X ]�L��<� �0^��vk����[�3��(���R��E��}^VCYi����c����N��I�(���`߬'eX�FB������m�sm��*��ݟ+�Cʃ��uSG����S��q���_�L{�����ڸ�["�ڤg�=½=��~�Ed���J�/i�ArT�_�Z34Dθ��:e��8w,ͬj�AN��p�_.�Q�㊾6q�,s9����}�>�
KOW��v C��*Ѫ�Z1"p�KK����Xz|v�����A(qݒ���T����o" ,����r�;���$$R�T��4� o��IxD�u�2�Um��ԗX+���������fP(S�)�e=�:�P�sqK��K��vO\*���#�k>�(�X X�h�?=|��O���\<��ת8����М��.�D��fV=CS����e[��e�ӡ�	���j���b��y��[�MD2V�^�����yS��-�R�V�oS�jD$���R������q�s��	�ԉ���:0.��b�\�OK�9�Z��ؖ��'�F�R���N4}�RtS�d�.tiGS����~��v�Jf��=s;��!Y/o[�����=�l���n�C7�W#V���U��Rn�l�W�+e���(1���2�ٕw9��"���V�V%1��!ʯԚ�k�A:�%j�g��J3w�@����a�5��ް1�2/�1���g�ʹ�.�KLKl�drKg1�`詸TL�D5�M��᫺��&D�&�m�g���뜀(���L�4QJ:;!���|�F��6k�d���IF閂H �'R�p��;�#ƪD�����6#7Z67��l68�y�\��F��Y[�~W��l�)<�V�9c��3}IL�w��R��� b^"pfs���Ȳ(�j~7��XѠ7OkRydP��F-����g��Z�	��<�K+_��s��av��3'6��X-���c&�ٺ�o����ς���������'��y�\�@h5��Gp.>����lO-W諴~	A.TMWπ9M��Q�yU
�%������N�+S�g�	��$s=FH@~���(+P5���8��|U���?�_*�0n�����8$�����-@��$��@S�����}�e��ˠD;ٴ턄-{�����1��M��GtK �U��%����h�
I�M�u�\d'���3Z*`C�܁T�j�%�&��܇��Yf���;�9.$oE����gR<-�}���b���W �c*(�rE�zH�r7�팍�"y�`��,���%/���I��:zv���r���?$2�6c���h�w��=
���~|'�'P�9<��]�.�O�}7�|}����̄�v"���Y�LO�J��i�����b��lL��۰�NH/�MH�GW�>�{#�G�| �;V��.��BqA��Ͳ.\��B�%9�����*f4�8�8�!3�V���p�ӧ��HHrkI�2������҂�NCۛ_w��xW6�$�3$v�ǩ��֤�bq�%!1ŽWw���Sc��� ��n�G�#veDl�縋��P��2�/ӝ*���EQ���TH *Q���C��
�XL���@QI35)�q��,���,v���C�:����Ͽ��܃��`����8p�+�tsm�f��b֦j�D�&lS��'K��MU�ޅ�rUWk�5m&��4��-9즾�oι�H�Lzh߮�E���K���CPVu�z�JG��F4�a����,q�����'�צX=�d�?�OvCY������8ֳ�6��e�~�n��A�����M���>��v���啊��SHy�Z�̈���C��!�g�KT�<%����(��I1Զ�o����˸!�4D�f�):0�(�b�*��W(C��9��f[5��J1�p�Q��Ыk���JZ��]�g2ޚF=�<���ް��4���Eڈ��'��7{��w�D�O~���x�M[��0�囩`�>�+��"�c>W�2�v�c�k��3�J��Y�� D���Q��  �ާĦ}��\��m6�`Ӽ�V^� �1�D�g�ȳȦ��+<x�(���N���W�gKR,0�d�멏���r�mP����q��.C�z�hX{3Q!R�Ik�-�<��`��Ξ�>W��5ڤ�:��˥+��U:���pħGj&;$�#^���I��^+Nr'�����Bu������o"X[x�h�iu�8̒b�eBu.�^I�k���?[h����J0�o:��h�:D;@�S �k�9�Ci5U^�D�ӻ����R�qɆ����ܽ7��\[��a��E�^<�Rj�.�u7pٌYV���mL?�z���aw�{J%Y��_��;?f�����@˧�+���uF1O����|�g!:-X���2ESr~a����.s1Ze�k�ͬuC�^�&l���+�^���Z�X]�<���D`�X^��ћbw��{�$s��9 M�xAD��~��(���)�QJ����o�
�Ǹ0����>d�E�W8�7M��#��2idq18�)�k��(��x������V: �0 4tC\�
e9R'�{I2X��"��𑠗.���"
1�a%���Lt�/P8���p�w��@N���n(ԍ��5�ڞ0�z���3	�$D�����4���Q��҃��o���w3kC�Ó����6S����jJF/�A�ɞF��=\K�Gn�G�"%�W^Gb���]<�W ���lP��F�zs��bi��e8V~��Jt��y(����p��l�t��+���Ѷ�_�k�IS&O�� �uȦ�I{��2�Nj��LS��+���W�q�\G�J��I��99�6�{�C79��&|����������/Q�9ċԂ�!Z)m�/K�xe�8Q�%��%ҺĹ�!Wx�ʴ�
8��J�=���%���h(K(��2,J�Z������\K��4���_},u/VV��!	�G�ͬ�����8] ��f�e(��P76d�Z' R[PҪ�D�X�J'�KA�\w*���+�\�@�l�\�SϻZ�/�8b;���Y���?�����,��(�R*K�6\�79�m�Glv$i!�����5�bȿ�(��GKD�{�UQ>�1Gl����<�z�"k'����i����p%NP���j���dL�RG���[�(�oXֳ�����`�6�>��V�l*m����D��J7��2�ye
X6:L	��J;=-�b��E�'����}�t�/M F����2��z�8'�Y1w5+�\����F�|G�N�"ҩB��f*�o ��P?�/�,;y@����Vڡx�V�.�]�ZY�G���^�#P�F�pL�$oI�;Mq� eɚ>6�s�跞���B?D����@\	����P��V�Bօ;&
��8|�T�?.r��o�j�m���4N�&��R��νHO� �
7��*X�lN=�
<���'�z�
�^��$w��Sˋ��D]ڼ��P��?�,Gm�;�0��-� ;��(<Ѩ�aL�J[���^��᫳*"z'�9am�.<i��l�o&x�;s@��{X-�6G,h�}w���d���Y�O�(D��fd��v-��1����!'}�P�ۂ�2W���s4�C+"PB��Y_�`i_"}Tv5I�@<���=J%��b^F`�R��dQr�Ĭ�U��^�5�r��]IW�S���v�I��{�� &��8����v�*cD��00� T(��X>@a3�v4#���KU�<��/u�����i4��"�3&��Dm���[i�g�ތ��G��3��i0
��7L�)�М���y�!��\��Z]i��b�����v׎��ܶ���C}X�:�^N�&3�@��uawyƅ�M�*��(w�]2��YTP$+��cΖ������\������]���	V@9t���eĿ���I%�RD!���>҃����?���V��>T���vT�R����0t���#��aj��X-b��8C��X�<W�}�n� A>+�Ysj��m�Uz��$ҡa�a����l��vh`з�����X�K���u�W6
&���y���M1x�.
�� (iQh8����D%i�lxi�L�n��6qy�n��^o�<�a�qA%	�
`�e~�����:�BN�K�NP4�����^�>�EӾR�ajL�s�����S4q�Bs�&�~�g��^�<�K�T���s�/�r�����aQ��0��3M�Y�^�e;��F��v[�^���Ox���q�s�l�}�4W�/�>0�p�d����2�@r���vO(4�
�|%�mdm\�;���Ck&�z��K�55�w��]�5�AP��`���7 ަ��E.�)y%Z����Q�Ʉ]oH�h%�D<3ŉU3��<O:��C�h���3�.aJw��z�s�����<٣DpLQ}���B�k٨���+W��������y�.� �q���<)�a+�y�dC�S#V�l8� �i��To9:N	l_���_�����4S� Q������1f��ex��%ۭ	��{�IXN/��1�q�"U�E�e��˚yc"�uZJ9'h��a���x3��۔�aG�L� ��ױբ�1�[Է;D���;*C��2�WUk-fM�#U��'��:H��w:�5��29���z�%�(����dSݦ��%�%z��n��� ���6�n�dufL�	�X�?gl�O��V3E?[������4/3��:<0,�l�ʞ�/�@�NP�I�-ul�L^��=dS�Z1�to"/��)����:G1��	&Yd?��bGA����8!z)
�Ue�8�%�9#��^��Qu���Q)����/~��	A!�DN�W�bk-.�[ΑX���j�&���h�E*Ќ�W��ѦG�ĵd�	���%B�D(�O�����r\�����I��%�K�RF�*�m��b��.,h�i��MJD
4�䎴V'�mp�=<b��wP�Jw����?�l1�ķ����3�?d�9kaT
	յ~P W�ɶ�ȓ d�� It������.I��3y&2"�v2�]g������M9�L��q�!=P��8bK��O.�����d�C^�o�60� ']�P��W�WI3ީҐ�mg ^��J��[�r�3ڽ��kd(��o|�$��}%F[�1��:'��^�$S:���}��@�^Y���������&�x桅��r�T��	mDI�J������nhiw��	���9ίJe�x��ퟺ��p^F6l�b��beS '�щ������?Y,�M�4���j��
00�v5�p1�����R�։�������ҥ���@�s�Tzi6�g��b��+���ήf��;��$-,�c*�޻,�]��v��%����B�h;�c��lp��ݗ t�z�R��k����Ab4Y��I	d_��^ﰱ���F�
�n���	�8������.!��g_I��\�Z���2� ���)Cwō�*\G�.)�ֻ��k���o�GF�D:Y��ը���Ȩ�BNm��Qye���)ۯ��U�P�%қ���u���-a�,�2J.�1�:��p�m�K萲�x��F\?|��L���j"����"��6Ľ7���皎��_��}[��t��M<ν$u�����ZnrHY�/=F�k"b{%QF�&\�y���Ɉt���+�a�^���"�@���כ���vX<�����<�����K;d�@�oY��<i�W((!��$���6��I"l�b�?��g��j1��\F�"��$~�#���O=K�5�ѽ%kV�iޟ��Y����z�ϫBE�jO|��$���X�S\OM6�^�Ĺ���?����r��4��_���RK�� OO3PB�d� �|m��~��#��#(IP���ܯq�FfB��'�l�cAf��)�_�9�2�Пi���6��YZ�@�g�������+�ӕwj�'�h�7\��;�3��Cv�+)f)��TBP	R���$ϭ2�t�MUV`�#�+	��)�T���/�ȹt.?,h�L�p�Z�A�L�'Dǝ�}c���+��j�*�w�DH�Z{R3�_�Tl��o���ʡ]Y_,�5E�~E,3�2���������n7W�Dw�/�0謾��"t,8B�S;��m�z�ys�M^)�5�E��M�4�/S��^<8a���pE�Z�֭.%�ac�;:�U�
���C�ZYH��Q�Rp�i^��H�1Z����֖.u���C�ˮ_Y�ב��f�+m<[���Ԇ��lk��u��K�$(��Ї�M�		�����Z��d�@2��W�TYt�W
FhxΘ�8�Ui��#����؎շZ���i�-�1D����sZ1ąm&46�g(�WkiWU��hA�N�}��x}��@���cD�����j~�].��vzL�5y�礪 ��Ǘ��H[ۀ�o�pFYG˶ėrn:^�lY&���Oj��?��!N�t�[��N����p��w�������K��]��D>�!��#jX�&���V!w�����\$�Tm���B�U�G��D�|q�k�C�j-J�%-m�W�#�k��~���H�_Q19�-�%Z9.0~�G�YQ��*8ME\��"����Q��b�C�I�q���+�Ͷkt:�ǿ���c	S��� �_���#�'�Y�B���Q<_�.IihƼZ:�i4O�E�-�-�okp��[A�/a���)~X���z�7����^�^{?����V`E2-�ۣ	�C�����,���ղв�#���+��� ����Mf�\��a�o�{�F9[Uir�4�Md�����A��*���\ӱ'FB�2�_�S�z��PF�&�O�������g8�L&��"T<���Ys��9�P$D���ANf���bk�Y��6�l�e�;�Qz+�Q;�4���@��0y��G�\V۠�JK����݉ɻ���Բr�&L{/R}K��b����T�ԕ��"�l���?2�N�>�(�������|�汉M0�D�\<���HF����*������C��'�y?�3�ѴQ�ho�㵁�n"J� ���W�����T��=�꙼��a�}�s��ى�e6���ӕ�$l����Nh&وF�fz����L%&k��6?�sgHg�	9˴��WE0�l����t��/=��A��i��n��y�dB��1i�(�9�����Fq�Z����zӾ���!W���w݆D�3nA�,�
�R�n��^��\k��t�1n2(�r-�����Roqy�R�gO�mk�!�N�Qn��n�ٳe�_�<�
5�T�������=P�'^��(k_�m�l�ƐU�� �
S��i\Yt���K�&�L�:v�/�B�4k��}��a������L��B�R׺�q�B���n�J��џrŠj]ؒ�k�g�r����*��ﶡڶ1��+\�@�����*�V��.A��f(E����f�BB�DA�{i	��f(	�zh�A�繾���̟9��^{����O��wt��И*�wT~���?%)ģ�<��m����o�&s�_p�:w��"���)����Uq�|��'�;����Lm;�ģg}��g�t������(��3�+�P̞����9IX�8���t�![��r���/BK���U̥B�0�!�����/�_�k���l�zVZ����=�Ŗ�NV�I퍊\Nò���H�,�;>{�(�������\�����˜S�?|9���ч���lR��lz|��TWd�'���SF��E��$�N�`��w�X�ٲ��h�ڼ������[G�o�U-���	���p����b&��	��������է��X���@YC86��o9�=rټV{�'%�Е���Gw��'V-ƃO%wU�z�c$�~��?Ir�4��>����<��&�:T� n��&�Y��~h�'m�ѡ�_����8n*7����B�ê����2w�E�J�3?���e6m��Ӈ��f�N�X��ֹ��~�a�p�:��%�<�%]�D2��gb�2���I�(�[�O�o-A�m���=������ܻ�2�2���UR��?��{�I�<b]f�43+|��2�@h	�q˽��uV�!k����2���G�+N�{i�I��s�w8	:T�Z�#���r@q4y�u+���Ƅߵ>�SWu��䌜�n����t�I�;�vX�U+�ǂv�q-�agQ�L9|O�c���_ͱ�t��Q��)����F�-1��U�ڴ<�s�$T^SO1�K���&Fu��&��6��|W�}�P2�D9{V��,�f���߇w�2�2�C*�p׳^w%���,���P sUw�.);���)j�4~�t��T@Xk���Fm��0�b�����S��q�3.�ذ�M䧅�%1���"���eݾ
�T�籇���n��_��ȚR!$h��xD�lZX�	t��7L�oӬ�:�>����U��������@�՚�x�=o����ۀA�f�ӌ��C,FZ�Le��?��["\V'��	��uS�3ȔI�RS����I�ՑO	}����ɑ���³�0����C�r�%C�Ig�-[p�˵��O��)�_����U�uݪ%��
��HT�Y96|g���Ǖl�����XR%���QhA�gL�T�$D�@T�MۍȊ���=DM6�~2���/�X�Y`ʊ��	��!w)΢�[1�u��NU��I/6_�қITY׈�8��ÚT��N�ea�u�ę/�����̀��$�sF���5�)���T6���w���#������z�z<R��#�*J��靸�ǜ�����|;�6��L�_Z�YL��@26̔կw��������S{(s�žT]��{���>�j���d��D�������/�u���p{+�)��w��jn���P�^���V�������<�M����
� ���]bskQ�4Ro����u��Y��A�aj���л�5�]∇�{�FB�+1_��pp�c�c'/,�+�o	&u��^���Yʻ@=��F0<Et��J��YYI��|c��S]K3o�:��	|��֎
���ur��X�9�D0�ԃ�K���-�/q���,-�A�z�6HA
�I ����$8K�� n�n�rleI��}��_,k��U��J"�6�х>��S�a��?�)��B=�J�zVNY��cf��5��v��3�b?��Cc#ļ0HqI��L�Y�vE�N����3���ݗR��uɁ�?j&��Q]T��,^�r���v|%�\�>�о�!z���7�*�%n�gn��|�'�J(�ɛ#2���#k�{i��$p�\�ȅ���X�@�T'����l��O霈��YڰJ)��H�bOBU|��^���d�<S�vZ�K �m�q�A��u�`����C{�s^��H���N".o���b�	���+y>2o!�٦��~C���Hl��K��:;�LU�Y�[��yg�귎�;DsPM�n��D���#/��/��ۍ��=.�����?�)3S�7�3I�����k�j�xP��W�}��i�;�#��{�]�D���+�Y$���6�GWa�z���
+�����z�Ё��߹ߊ�X���_�ˌ�����f��UT҉5;T��f?RmJi�kx��/@d�r��Z�"r�z�)�U�Q�o���M_O�޲�Gk��8�^���q�C��.`oeŗ	�R3A�%'̫��d�IU�����[���ɚ���S�A�9l1*÷�Ҋ8ف�{tf���*���n���q~�:k���

H���4�&i�4�׭�~�5��-�z���.���60�'������w�45B�
�n��C{	 ���������So8��n���e9��������O�5և�ǣ3ر��7�����[��	��K���;�*�q5	�\z�j
�3��R�8��Wh]DzM�����"���8Lc�����@U����^,C:,8���$��N��*)G�j�.�4|v� �N-?�r��5r��l���[M@�E�'{[��ɾ�U�@�G��8����E���G��8���G��YQQ�� ܛB
M�/�d��V
���=d�%?
jYw|AQ�->�R��ƏU����^�Y��g|��Σx܌Zޭ�и�؟+�t@�K������m�Z|�]�
��H)����:�\�B��������v�]\k�����iʆ���-�:.kT��YX�m��*��0g���$M����2�T+��S^�&���w@��L���K9��bV��w_�j�AthH��
��uȨ/?S�S�������Ϭo�ǃsk��(�1�-�X�:�p�4/��9�<?�R�j�AD����`yS,˘}���8:����%��>���(�#�fV��).�������nN�8-D�$܏O��H����+���E4��>"�5���0V�|�r����/ٲֹ��+���a�IE98#Ut]�f�2ܣ,�ʻ��ړ)����5����0�����`*2_�`7C�]m<e���F�µ��}�p� T�y�O�1U��:ݑp?�[�_e���{�շ��M�}m<"�NG�>��I��6\�c��� �
�]r� ��e�����iE�Ʀ�gJUiEnj��R��0?��  ��ef������jK���I��#$������p� ;��X~&@8˜�1#J�fMÀȱ�V�t��	��(g�XY#����7�g�E�9ծֲ�Ψ&�����=�u̲��SNK��Y��Eɸ���R���+��M�c�z�,}�zY�W�Cy->�l�Ya��AK��"O�̦8U���X�>�Qm�%�m�<� �x�?H�]f�3O ��d��hr� Ex�]��*��Ƃr�Q�۹+ �K1�'��&=K&6���l�O!����������]��]��s't�<\�5���q�^EXҖ�)���<⧼ �	T���~��.: �q�I����S�C�ڊ�_Ǽ��ʆ�ѓ7�ZsT�'�.�3	��	�&E�rE�o�nfPl��5�c��uVz��(kR�W�t��ɡm�qIx|�q	�������=x����5D�~ sAiU��b����Q��JC��J�[f�ZAx���|�	�+$l�dW�/f�����!.��5��ˎ�~�W�0����6[/>�]�{d�7]Q}l�ܺ�1����{��Զ�Z�ﭻZ9�yAݾ�F-0������!���:����t�oZ8����������Fi4L��~��:a���Jv/�Ip��UEҌ��;�7kگ�B��m�=mV����Z����k36��W�	oXg��i��?��%�b�
�i�bf�t�1h�C����ަ�uܳ�������ț� ?ǲzV�o\eǩ���ٛ䀠��:~~�����k�&=8B���E�ԩ�=K�SwUJ{��7
=:�������5M���I˛ym~�w���f
;̬W�l��}8$-Z����N=����?秘�Y����V���_'j��C��8����ZM5���#}��z��oa�r�W<�r3<<�����eHxp�8�>:�o����z�^F�7��E��}�2bbb[����V�����m��~��G�}�":�^��թ�杪��"HZ�4V�4��'>����n;L����:����!55�]�M����:eK�szr��;��B��a�a�m�O�@HC�]��0��b�����O��4��L�)I�[k�;����qDh��pD�Tk�_�ߴ�J�,ڊ%������rd�{��pf���z�
"��5�&o �AS�/bߘ=㖙b~���bs�`�6w�i;fi����(���߽u0+xC��
}��Q�a�R�J84+��A��.<���z1��c�ώ�>��Q�x�<|�a^#�h��6�w,���y��@#��yF,~�<�QʿL]�?a��c�;и71���"�20Z�K ł/�q��,}�W���Xh�{��?	�*(X�Zp��so��#wN���ޤk�)\�!$inl|ӝ�o�����`�ֳ@/��y�>�q�'�������݈�O|���	�4�<�X�A�u	p�"���O�x���k��1 �)#0�{��a$�z���e�U���D�,)ÿ�2z������)Q���7�"�?����f��\���>�ٞ�^�sQY�>���ӕk�]���R[M�a��WNT1��$0�U/qF��8ٰ�.��b�HA�A��_�jVv���<n,czP/µ�����(K�s�/�����V'�P�nڋ|��}<F֞�ڵ���og�P޶K�g$Yo����6,.U�w����	h�pcf�ψ��,���I�b�_�>m����ʻg�PC3O����7�{,c'c/�MbSa���ċ6��{c���Ɔ�Y+%�"�i}iR�X�z[yŻƟ���a>��)�iD���9�^w�[�8QIg�ŧ'F��Ws��Y��],�bB�cHF��b��/���|M��g�S�Svs��M:n&* �7��t˱��fS|���~LQtho�Y`Q$!����a�2YN��'�(v/"]-��]�0nW���_��b�@ب�����*��"�zNuU�մ�g`��:6�7���'U%����م~�zP�[voG�x�l�_�U��R3=��� '�ki�1%�Y����:rꋾ'��}8�	ˊ;��шE���Pس?���7��3x���I���>���y���tQ��"��K� ~�.1��4���5J���?��³����J�`$lvil���"B�ǳ�Om�-b��ʁ�ZIY���y���Vn�����i��;o;��=�z�t��u�d;6�I�-zj����M�݁�@�7�<A�^����o�E�U��baY���#_Bmj}S�R���u��Z6����7NW���z���b2k��B^M�����_�k�PP�A�Db|�19�A\�E��J�n�Ix�W4�/>C~�-	9�_�Jɔ�X�B�MѸ�=+�����t�u�������z���4�-�{p�ML���G�,'Ye����[��K��|�$�={Z��%�ny��hY����R2?K\r@�7U�����E��ƐE���
�t|q�����p���O�*z���0��z�Tt���@X��%��'rߤ;��[��5�y���^���=������l3�W���5�̓_�8�w6��/C$�yE����;k,BX��e�|��0�X<�T|�>�?�	�x��I�Q%���7j8���|�m��K��5������c��WG;VY�AIͥ��j�Lש�q��,3iM�SA�a^#��R�UJ_�4Q���7��K�b\�Oc���>L�����g���'(�H5f���W�)d�߄�w�ȵ��7�Z��B������f��0��`4�ܕ������;�([U�=��<�1����l���3]���g{�5�F�i���oթ���g<N��X��P�%���.���A��b��hвq�,���?��Ԭw�j���n5�ԑ�+�\�>?����|�u�t�J����U��G}.�N� `yZ��O�Q��~S�}�g��dF��`�4�Eg��Z��Iډ,�,�U*� ͫ<5X�A4P��>|) �|���>/����R~d�eDC��@ͬ{(�
�>�ZT�.º֞��-.��ao�m@3�����0��X�@w�7Ҭ���`���5:�y�N^"f̼�V���Xȹ���p�[���x������΋-!#wa�e}���]�>�z�iÐ�N�n��1�t��"%��~��u�wb�̫���r��5�7�Z���Q(����%CCjum�����Z�h9	��AGR�Whp��u�2�8B|γb�o<���,��7y�0�� �a 4�d')�;�u�J�����r�[���8�v�Ƙ�l&���=L�R��!#Ѡ��O���Gm�ҺN�����%L��Z�RoYo��r�\����(U��kk���Q0��=4Vv��D�U��0/�!RN>3NJY�h�2-]���i�����W��0V�<�a����7j5��&"��R��j�)��s6��=��~{9����8R�A���e�ݘ��Le�N���0�C��&D4۟:���e�D�ay��Dk)(�X�gj*�Vz�ů�f�t(/~#8j��C�'�E	)��2�M+�ҭ��x��z������֣;�����*�H�V�J���4�~ 渘����w��9����R��h���Z�F��&,cdc;
��Pl��2��\H=�#��i�A�`~/ ��s�|����Se=w������v����[�J�.�č�}HI�tKj��Z����2I�p��ZvW�TN]�n�Ā����/�̛9m�؉D�XՔL9�<�o�0���:uN�}�U7�i���',Pl�_MM,SU��)Z����y@��\��/����"y�-���(���y�P�~́yu� �R<�ԀO@�u�a9沦#��Td>��{ݳST�8����>/�S/,�>ƫ�"���٘!�4��
��4���p��>En�bP�B,�у=��g|�*�9ۋ��&��/�B:����:m|�C2d���l��i9؍��	G���_�<���b��փ����1���i�P��%�ǥs��;�q�M��*�K�4�5�֒ͺZ�Cɻ�}�����Y=u��8{g4�)��~�e�mVf�g��Ҙ�Uf�(��}h�^R)�����M&G�$��m����=�ܨ�{��bT�O&�w���t�ޫ���!��÷3[�X9����E� 2��z4�s���.7��4?o��+o&�7*�8dF��+c?��I�}���A.u��p���������{�?8�È���疠?�7��f{<W���9�5��*b�i�WQ�������o�!K�V����`��
x����G0������vd���楶b"J��]���J26�A92½���C7����n6�d6Ms��)@ZK$C�ᕈ^��5�w"γi��ח�1x7_ '�ZOa�y�}+3�!���7v��r�	���=�$e���e}l=$�?�Y�����\�=��l���zf_��*b-�6�Q��q�Ѻ�n�9�2b���Lc����礓
W�F�c�$�9l�
u|�.��]R{��q|W"/)���}���.T	ٳ��#�T\��1x�4='��w�AG:{'RW-Z@�v +�j5����x���2��l��e��Y�; �bnrHu�Uv���i�
��<v;;;s���18�M2;�[�{|��2%/�U�C���-�
H��f�.�M�'.8WE�uQ7��o��2C9��gIm�~|kj�԰I�hg�75�Yyxŗ�c�*g�nw��}�9m���Y����83OXG��008� �푴A���~PY�C=�u�����_�#5�yp�}�I�� ��w ��O{�����r�_��!�hʯ�l�-����qoڪHp�"zt�̴�6Mr�e�D���2J�I�	�N����j?*���� (����a��?/�d�$�3g�02�Z��b��?��mJq�}����^����#��c2��P�h�u�qq����oE��a���W"j���ǑI��-U��K�[��O��	�ond�O�&29F	�w'ܴ
�%#�+�^���ӜIi��Ȟg�~�f	��M�T�~뗩��{ g�I>�@-�B�X�߀���o�ا�븿�n?�0L`����yϠ!���q�,P될q���3Q �����F�p߈қdK��.xNA���U�aY�Ӊ�7��w�䯫C�����i
��� u&!+�1�i�F��k�Mv �[�:�IbTT������$���ƧjV%����s��aJ��0ޢ��T��"�X�J����]�k���ˑ��b��+��=j-�,;m3���-#��[�*BS�4E�L��J�n=?��p�l�����o�����p�^d�j��
ӏ�b+kk>��'9�;�
8T	��~���2�-wT���46�p�y��4�ֆa�U�6>Rs� ��y�L���F�K��}TF�c��*��$4�_���s5m]���R��c
�>�E��: �J!�:���t�2���4�.�[��mlX�.�giߞ=-G1���6�-�U�Zco/K�+�o2H%2d���u���}����eӥ�i�%���e�H�U�<m�Ư��S��ъJ�f�ce^�?��8��t^��p��0���n$�}`ո�ʣ�T�5 Bd��:�ף���
�{7y�i'��@u��)��X�	�Z�u{�й���F�ۆ����ޡ�̿6�1X�k�KH�JH�N]�<VId~�
�
�2VϾ[�h�?��g򑼅�{yF�L��D�'d`iŀ[M�n&G�#k)�e�K������f�/��=�=�d���3��>�%X����
~f晋]�ӊҲGS����~A�H���<1�I� A����������BDB��k��%*���]Լ�[7�Q��X�i ��whi�g������g�0�C���"��]�f���2���*>ˇߌ�y��.I�T��f,�U����Oߎ�Z�W1�06�\n(e��셔R��du��1N�嶫���h���G}��X��w��q�����~�l��� {���l�5[��ہDv�Az�OnZ�f���;��W�
D���ׯ�"�2O��)~*��3�U@���|����KK��I��È��
lʫ� ��	�S��h�+�Q�X�h���$!A��&� 0��3��vY���=rN:����u+:*wY�����Q�~�I�KxE�EdݑN�ܯ���>!������#�+�q����&��oԹ�T/��1�w�����_�Ft�D^����2Y�����6�9j����%hRH	Rތh��A�/�`ۛ�ra��ZG�����=г��ExM<�y��=\����؇��%�$��w�N��d�u���ۄ{PN��b���+����Ne���
�x�{��r����}]���Ayd��?�sh�������L�\1�yL��[Sz�G��&=`���׸t,;��fɄ-�M���۩<�K�^�#Veggۉ����o��#��u��S�S�B���� 0|�W�#�ۗ���~�&�+*$��ZLj9�:4�8�!G�T�S��7ٟmB&�L
�Ǆ��8���M���RE����}]�R�lW�߮<+>"�>�yX�yd!��X���
?�c�������s�e�R��rX��Q�s��9��3w��)�E&�aQqp?���� �5#omMG4���E+���%�?D��x&0}M�d?�h6G9��
�I��%'2�j$0aHj����W�t�ϓ��0���:!|���Ԕ*Y��g>h5?�̦���Ŧ'
�:Q�εg'�"�_�,0�[�@��\>\v=�,ϑcǅ@�chB��a&X	���O�]>Թ�QK˸*V�c)Z{4�-ځ�?b�m����6���tE�BD$)�_
�hmOMi�H�1���7^�+@��Ƣ���'+yv[���$�_^�&Z���n�ݑ;/B%`�%��}��UZ��ZN��k��k�Є!k�u������Ac�9�z;EÚXD]� �}�͢����Ï����GD>��]<���-f���m(�-�)o��?��t�����C���|�34O}K23^��D�;&b�v���T��E�M�����Nf��D"�K�o�-�;k���F5C^��蠲N�2�^�8�U�H6�f�����y0K���ڰ
/թMG܁�z��&����[���d[����)����.�6Vb���AxG��YKl�W~��wH5 6��h�D�L��jV>=��( ,�z��o�MR�`i�Y�[����ad��j�HS���M2b��[�xg����Y����3)F�t����eN�ZK�%�~ �w3v�eC��?�ʞ��&�\^O؇�x�r�:X��XK��u��a���3������[ʀ �jM��K�q��F+D����|iAQn㡲�ڽw�����ɓ#�1�/Mg�O<�;Ӟ��36�c���#�߻~��_��k�s�y�ʶ7~��L��u�w�T���Tt���s��%:�Q�M=��=���Ԏ�Q�H�9��� �'�\Ȣ���Q�p@���� �_o�H�n�/"b����v��*�5��>�f��S�k�V��y�:�W-�R��_�AY��qxxxZ�(�Q�Ry�������A^�����
G�[����73�3�#���7���N�5!j�z�r�󧟣�\ K�^�eo,ӼsЙ����3R�|j��j> �uW����N�`r�+s�*�Pur���#��*1�h�]��+ a;@ݝ����7�8��h�!d'�E�@\���l���On`��^>��K�42D�z��=T 3���l·">,&�Z����&b����a�#���o��J�ť�d�\J2Uq�f��jL��3-���Xz�Q��2�[��<�C�Y����Σ�*z����ۓJ11~/1�ꌛ�r�Z� Ֆhf��*4e�h�P��Ɓu�/��C�f�B�?��o���Z|� �m��M�^��)�7ɗWuum��~9���˻��֡��vl�<l[��$�S�e�+ü4�z�ś2颕�^l�.� �U�
*C��g�9:��jh��yB_��;(����7�CP��M(s*��;� �5���L`}ZќM��|��[��4�
�����* ����_�i���/�ͯ�ٺ�a��o�~[g�(�dP��Ö��m���6�0���xc��_e�Z���|��ј��C��X�4�FJƄ�:I���S[�\�z�˝�_�����}UqAՇTtF�V�l�AF�;(V���4�uǒWP�b&�&ɡ��c�V�4����{�� m3H�VW��*�ÂR�z���VX��� ��k��׊&=�"�|4r��ׇӏ:���3�$,�N�@���#e�����W��y�s������Ҝ���q�0��<%epz���+�߈]D�\�OqU�X��3��a�QE>�+���ER}�J��9���R��B��G����c0���b|�GqV�z��]�X.�0��8��Z���U�1�o��+�˃�i��ʷ��@�����Y�㖐�o,ٰ�_"����<ǣ���*�M���,��i��	EqQ�H@WH����{X��ƓO����P�U�uum֡�ݝw� *+I��9Ľ/��A���I���i��s�v�G����Ɇ���_y���.�x�9t��\�#BV�|I��R2�������!/�7�j��G����ΠoL���������8�:�%�4 ���LH�۴��SDM,���+5ni�-��8����/(A��5����,f�3ʤ�ʪ�v�����p-��喱Yl�?��X�C�;sV���N������l�] \���&أ {(��s��j�Z�ϴYzݠ���CV�D`.�Ğ��'��8��}������$�c+�F���~�����~סwU�F�w�iC��\>Eq Qד�9+��}Yh%3�/�U��^Y�Pr'�������c��:�;*�\�0n��@�d�'�t���++b}]�?J���[���j��(YԄ���k[�w���E���%H����I~��/�������ͺ숙~�d�﨏��L�d�%6%��/�*d1'u.9�|�aFS�����)��YA����d�? ���>W�)E����t��x�~?ow���#ɳ�VÊa�`��B�������>��6�9$I;������?�뮭�����Le%wq`J�~�d�E�v�-��JN>0>�Y�W�r�[��X�~O����"����l�5#G�83k�{
�Ӣܛf�%L�?q�|����~���)<T�N�J��PG��Ki3�����!�/� �[���D3ؖ#�}HL�3�᛽X�����Q[�n_|��O��!�>�v�9�ilSb�����@��y�-fI�33l�wG�;�j�����s�?6��;�bV1��#���y(ՇRfU+LJ'^"�B��vk������B�	�$x1�uy(j�`����nce�m���a�Cf��l�ڿ���2vӠ��Zm7Z��H_qZ�P���د���3$�v.���.�SU����;�ĐrD$}cٷ&P���y*x�Lw!��rlHL��a�8��>�tM;V��͍��D��W�c'ݙ�<)�>N�jk*���%G�8�4��wR��w	l!���`dR�AW��$ʿ-&��f����2B�������o��.�����_uG���o`YC�M5=��$�z�H�.bS�sC��e��/�Ї�Q��+��+�wD����l�k����'0��C���\!��P�)v�{Һ��u�S���,�>F���}�B�� 륧k�$B +�-E������>�j�A����>Þ��a[~�����ǅ�����]s��~�5�3�UpY�xw�6�	M]o>rh�kV���:w����pu�l���Hxe"oؗe1%��P'U~��4� �
��g*�&���c��3�b%`O3��'��y~��TOl5{3���wm�s񀟯$d��*���6��*��Dx@UW�*�P}�5<�)[��1����Ow��u�]�LH8ӝ��!j�%�_��ܗ�2�`՝���tԀiv]�C6%d�K�Շ�H��zt�w���Q����7�e^�.^[\d�пEZ5�<j�����IV)�ʊ�����$�<D�-��_lB��/3{��"�0��bp"ry2+��A'���K\� �jNy��:�H+:��蔳EQ�[���T��q�n1s��rx3�\��W���o���R3`��^�~r�O��5�j�H���Wj��w_����?t{0Jh�A��+Xh��L��`1}j	��5z���'�A���#�c�d*� 'A�\�f���#b���JKP���Z��9�վ���'Z�^�/.�98�r^md������2�x�.�n�φ�������YG�G�������'�)@9�����/�@)洆�D�)*�CB<��O�d��H���	�5��ʀR'|��uZ�%^q�W��N�X��n�ⅨXt/Cg�bݢVp�[Y^t�+m�A U����1MF��&O�3��-R��Ӽt7����d�4��aZ]���U�Ȧ�B�c���{�Veo�a�H��J\ȣ����oRk��s%e�[qi�%|'�;+�3_rX�
"vGNW���|��7&%���ߤ��k=11����m��:#�������?ox�+8�/}�c�}ߒ�튉����\�*��A힇چ�s�033HW�?�%F�UZ�k��R2�t����CC�({e������e	 �}�s�Gwj�S�f<�ƭ�$~��O��]��J���B�"�ɷW�O�ϮAM��i"�sv���"�yS,��=r��s,�L{�5,*� �p�  �L^8�ԓ���,B����*_�7�4��/�3����42M|���8�8'�+9�6�%�λ�/�z�k`�7���]��J;|�S�5���A�m���������u��iR��,P�&��zR*�%"���B�kfjI[����c�'����B���<A�T�°��${ǩ#s��ܞG���3�U����1w�L�x�\��B5"�mV/G�]^�z�2����o��|�g�����si����?��z^{�B�%z��]5�+��/�iXZ�T4H&�ht���ڣ |�Y��x���,���0PG;���0r��i��2�^��l��x�Jv+�O��N)����T���<��FP`��%�o�!��&���Am��ky�%�߻l+�8H�l�
�/��Uz@c,�ư5!�8���52ɣ�����UEX��ӷ9�˭�,��M p~�4i+tకU�-]#�l)�GYQG7���Uo�>}Q 5��M9�B<�J�0�d�w�8��Ȩp4�:`x�:��j#���^�A�5��Zxe�IďjM��s�ƹ�=����x�1C���"j��dk�oӆ�j��S�������^����l?��-5B�yW����KG�5)R��r�`��XxAԜ���	�����wrN? ��YI2�����L3[�r6��V�u�?^��A�a-���R)i{2pS���f���~D�~%���
��(?V�s���wS+�����_vU���c���T.)W�q��`
)��oը���ϯA��s|�Dt
AU����%@E�J�,���U�^��39�t�HT����v��<��<؝>TD��-輄�m}��Lu=+�]�l��T�
�ɡL$�u)#EZ֎*&a ��� ���?��&�'��X���D���g�j�%��o��	_%J����D667� �� �];�=��ڜ
����/���E��VÞ�y��i���~��	�u��MлFz����W�4O�.O���eӬJ���9��b{�/hxfh��)����wp =s��c��Q���n�v�a'��)!L!����ϗ�,���Pwi��6_�dD�)�5 ?����p�X��b�R��|���!q3`o�ޅ����� ��]P������ya�X�p ������SI����u)|�c_�(�7�#������O���
��zz��(���P5(�X1�.�bU$¡'T�-�;�FE2ь�NM�$���>�UV�w"��[<s}���d�=��rW����޽�Ks��V��D��{ܕ{7�h" �ń���{%���^�r�i��>���0�Hr�JM�(�[4�\<��'�-=���=�&��h��l��aLs"���?�k��~1 z����m�*l�a1���?�醙=���n�N[�k�Y�e�"�x�U2~���O������A,��G���x;��nU�����Z��˝�峒��)�e%�l1Zܛ�Ȁ���i~7I�T�2�z7"�-� ���C�
��_蕼_�����0hU��jv�� �������g�t�Ǥ#P��󿷋(dǌ�\��rU_�P�J:�qD����'�<��H�U���%�]�TUN�`='�T� �=��0�
�K���c��6e��Q��'�N�+�J�!�c~����/�1�rd،p^���"��&�i��pcƐ�ꧡ���K􈾟=��{�@�`�Z���N��,x��������p��%������̻wr��ܹZQ����� �f��aU�K��jcL3@�̟, �U0��L�k���>�YĆgTH�w����*K�p�n�=�4$E��P�㷺l[UxFtlp 8WA���Y��-��g<e��yNd����$k��Y�ӈ𻆉�(��͡|�����v���"��ѽf������
���'ݖ[�'�I/�oз��wV�s�0��u�k�ul=Z�r�u̒���	�K�O������{�z������m޻�,���j^/���3�<�}�Y�OC�ugm�A*D3�8����q�c*kz�Я��V��r���lR�{�k���/�sa�+6�t��8ӎ���ƔR=o���o�)�0W'��q�!��<�ז�-�8�,�����;�|��P�l�g��K�❱�1]h�4ԻP�yK����>�[��/3�������Mw��I�l�D�>s������mp�޳�59������r]5uuKGG�TU���|>T�U2��ꢟ>�Ud�2Φ�����Z��l�
=�K��T�4�Э�p���x8T�w�b�&���D�\��4#B]8�Ӧ%��y�A�s5.i�n&�>mU'���5��j���'ٓ>[���j��C�{\�d���a�����#��N^AW�nvv�:��Ƥ�ώp�Ʉ�s�V\�櫛�\ѹ�w�[���_s;���Ͷ�����!��N��W�P��eb H��R�K�dd�.�T�ȕ6�Ȗjk���ՙr]z���;u��r�	�&`6��s���ɔ+Gz9?�oc���L�h6��5�W�iu���1�t�Q�:2��'��:s��>��a���r+��9�OBU�n�t��m�,����9[^.�5X��e"I���)5�;��[s=b�g�\�M��L`'��ʚ�bᜂ�~�c'-��Q#M���Cb��el���?G-y�a�E��������'^����QQv�ޤtJ���t# ) � !�"%� Ҩt
HH#��J#��H3C����u�\�,������>g����~�����w��qț����Q;����kO����[�$oo�������K���"�|K�= �$}�52%�nw���;����eec���UϜ�0�;���0�7۵�����A�����,��MT��~��"MJ�Ŵ�ʮ���S7Ѯ��9�˲)Ͽ�l"���#�:����aò�sM��fb�����ô����Pl>~��S8���63H���	������6/�:��S{v�EJZ�.o,Yf��i�#`'��|�QG$J�J�'Xc��\��d5��#���) ��K����Ff>��}� �Jz�7�X3�Gk9[�"_س�E>f��Ń����]f��𴴴\dZ�Vs܏���n>~l��,��a� ���ii���%��@��̖Z���xD�R����*"f�r�b}�-R�8��}��Q�(s�!9�)�۽��ז�8
�Ƣ��.�E��A�������>�2-H`-G�tF��($���w�|Q�tGw��+a�S޳�P˭NP������hL���Ԣ�� ��Ym�Qm4�	&))��������e�qV������#���^���с�Ч �gnVu7��ƫv�O:T)c�Q�n@,��\�fJ�H=<<$A�ÙOC�i���J���g�F���fJ�ah����u&~��x%&_���}d������s�ǣ��e���n�<Z�C�]�<��c�rE��褁��V̧�Q���pU�i��3ㅯ�$��4t�G��� /��uyN��eL�f���6"�OMuup�f�c�K��(d��<OcZ�Dٿt�44;�ҠW�/)�̄3o��T����T�^W��2q���Z�tKv��6�՗s��f}b�@i~pr�����rfaNk�]�f ��2j7ˢ�C|n�+�J%�/�4�e"�+4��-�%Pn�ʆ��7���^;T�jO�trf!_7��q��I�s`�m���ULrQ���|j�Z?F�+�0�-����+��u���[�'�9���?g�m`X�O~���z�9�w����܁9]�����s�*Sh��U���|�s�D6�)1��b�[+��>Z��b7��k5����X�9��o��k�eh���0��Pk�?��D&ઑ�$��ۡ�!�S�mmquuO<�lV��D"�ūm��UU�Oͧ� |Y�#��o�t]�F�ܛ����L���_ m����o��j1F<���+yLo��Jj�'h�_��ԧ����3z��7H�$�F?�]����^<�D=+s��'l��w��(¶S ��"��5��ȡOG$���x�@ȯ`�����>�%_��)O��c��4k�D���I�(U>�
잕�;���X��,�N˿�Z�)&��cҍY?�.P�g+���Cͻ���d����_SO/|��n�c?�tuu��^����>h6���Ԅ��ޡ��u>�WCS3��sn�=�A�Y�Q�^�-^�3vK�����@�Ufʂil�3;�����9�^V�:�N��B�}8��YT>i'��怲��A�!E�x�-&F2�f02�e�/x�
<�7��c�#���u�1�����;���>�Pbt=� �� zSXD�
�1�/��X����67�.\������nF��(��<��HWF��]��ߠ{�3a��@� 􀞞��x�bjj���9�/�y��@�nY�g�St�C�`�@jNN_��4:gL��莎�]W�*L�ြħ_>�)��`~�jÇx�9�����_S��wV�J��d�AZ7��ٞ�*���~���9��b��Kk<���q��M;��(�b��%4Z+�mt��ay�ƶ�gE�������5�N<#r*@�T��.�\1*hZ�L��UiZ>�DYZ.E�l� nĽ��M[�oib�e�ep�,�%�7��[�����M���d|q��_  <<L�-�Z��@7&��� +,Je��g367ﻸ��%�>n����Y�' iMZ|(6GrPp��GF�M"����t��]��h�g����HI���h���:Z#hF����A�G,hAY��/ "�(����f���lŵ�g����׋1�x�,��p^�%�E" ޘ{h_V�;П~k��SnI�F�O��A桄 q�v�n�+8�nL���|�飈�>��w�]u虁�3������66��L�y˞݀&605���q�����z=�1l�A>B��T��1]a�Un��z��O��F�-���#�S6Dx�����W*OВ�2YŃuٖ!b3V5*;�H�}��X?��4�����~�F�ֺ�8d�����}�S��c�ZksZ���<'ǳ.j�l'��˝�J�S���������>�r{��c������^*��r�g��ֺO�6���}"]A���3O���D�f�̓�`�吻^+}�;Nd#:Q!~�h^mF�o{J�k`h�17��I�#]c�/}�X�G)����)��?��]Ox*���x�+�C)��{{{��2�T�"�U�b�S��`�Xꅗ��\̧�;MJ�j�=�o�}>��J�1�_��{�>��*�<pd�,�e���a叝��|��$~U˿���� 	~�����b������`��қpo��^�B��%T��`�=�!"��Oaܟ%��9���Qr�|ի���ᡈ��>�7��m %hii���-'-����X��ֲ$i��o�f�rC�u�K���Zo,}�����|c��t���� ��F��CEQ�FɽI���ū����l��?�y�Z;-CstAA��ј��7Y�Zw�Ozo@��ˣ��C�J�ls~N�ƚ55�2��~��C�rys����;z���@�O�(�ڐ�� r���đ�;�E�9��Z��&i�o��Cȿ������#\gD��a���������r���wAe�k?sO�M���F���1A�t����,�JMH���Nhe���/%��Á�����ttt��<�4n'V�����Gypx8o�é�M��+�N\�z�<6C�J{,����N�A�rV�
�ɓ7y7�Ƙ8	>��*��x/SD����Ҩ�9����$Zܺ���AOi�$����=`�Vf̀Q&E��:7%H^#s���� (X���M�8Qա�;�ڢ����v;��/N����^�&f  �tG����4r�t�����f`b�`j��'���P<����s��t��7s�Е��K�r�I��vO��oZF�LUܲ�c����l$^��_nk�9l�nT,py�:�ȥ{ѝ0����\+ڨ�
p�n�~|i ��hG�e��Q��y�=��WeQ�L���g���۳?~J��}�nnL)��w]�����%�������K��P�w~/�Q�E�cZ�R5��+����^6�{�ō���~h�������$Wpct����Oԛ�����f �	O�1ȀO���� ����INIA� �D7����(n�ۘ�r`�%������H�p��Wfw����i3�+i[�7V8K���F��_�џr����h=�v���	t�l	8�ep�K��COXxE�O�G��m�;a=�@2��F���uV% �~�[��%ߗ>���c=�`VL�2���)���:��R@�A���%�γI��P�/�^>MA�#����m�*����p�V/�}ח(�?�9ܢ�����H��@�q�L)/B��cJ��0t至�}��S���w�s��v�PN��p�q�*X���=t�2�8K��l�Y��H��|���^�^D=�gߓ�����[w�ۥ:��";e���Z�k��j���K��5�z�T�f���N2~gBcsJj]�Oh� T)M�����_pnb\���-ݭ��L��y9�_̅DD��RgȖ��(U�I��9��?�)#7�aNh�$���Q'j)p����Kv{7���R4�E0�[h��<?����:�Y	�u=���voڃ�`�E��������^��MlΣ�~�]��}BV����"��~#�I��%�U��6E�#�s;�q52ɳ���yG��`E�N�����I3.��Rh��8����ӿ��j�u�B���G�<[˷,�z�<���b�;ńz�6����ɴ��2f�徴�ѐ����L�&	���M�s�g(�����bk4��ň�����m����h9aǉ`T��bum^�*���XX�2jE��C�,j�S}8x�z��NAꣃ��W+�?:ۦCͱcIb[M[D[�����&5��j^����|�Y����7���	����򙥚�������b����b+���?���i�d�>��������>\����*��4����1��/ƃ��]s����\�1�����O� 	neoO@DDtv
sAF�_a���S���ښ߲�����Kk ���םD���_O�]��kQcHB�������o��\�>�]�uchb�6v9�r�=���`gh;lv!�Ȟ�i���������.�M�,!M��j$�"��;��l��j��^m�r�v��W�/뙮�����S<i�@���O:9�ϾȪ���Y��6?�9Io��u<ʬ4;���<��I����� �c'��ߗ%���o�<�n�71�ۥ53%���A��pX���ry��xԫ�]���4	{,]W���'�ª6�L��ʼ�
�^�����5���0�@]�87���Ah�ǁHP��5���M:���y�(�v�m(_�.��I-���gE��6�2���w����MЋ��vpg�>4)}����i�MK�S��fg�ox�+��kvN���>�D�ܙ���E��:�����3�U����w|p�S�l�8�7,��\��)�uF�?)DHOQ��N��((���oֱ !��	� ��l�To*���$�ഽ��v��7��-���=Q��Z1�����P��}ޞ���$�Dm�ry���8n�\�Ϣ?��%���{�������Sy��"��*��Ȍ9l�%>=�t�<c ���\ox��:�������S�r+ƪ�>,�zB���g�.G�ss}yvs��4����O�a�ێ6l������4�z�T��>48��oӢ/�옂�`�~��<yA���`�mgC5�;! %!	h����X�G���}�� &G������������e.6lm(-��dI�������^�0��c����uO����tbYe%��.�ٿY�u�N JK���f{d&��!ٹ?A�Tvd{X�_f�M�������/��6��cjhW�||#�)#���`o��-����V3"�55��)���hU�Ԩ�fF�cnݐ�MG�Ю����V�ǩ���?>�=�yJ���5Ɔ.dd@P'Mz�#/3�s�;�������W���=��3��%	b3QOڭOV|��4�^dț�i�"�q�,�������Ht�1Q�y^�M@]ԏ�����M�IK�E���=�M'<�<�	�~Zi����1�gs�L*��� B~ڍ�d���#QMMM��.����=neee��b�;�+�-��5���OK��Ùە
��W����hB�>CJ�wW��
���-�t3]�	������Q�zf���{LWm���ee��}t��}p��'9^�����@�W���N~��g(Dk�j�]�����]��W-7�,��⻊=Z<�����떖������E~�������#������c�LXO���� 0us����=�~KUU���5`7�I�T�rc����;��y��&���m��w������R ���Xy�G#�(��ió4�A���c���x�f1��Q�tKU�^䞴IVM�7� әL���1�K��ǺW�Y=����wa��G�e�I�ʪ�Q�sjm�vn��:uD����I�O1qh�p30�Y\��)C�! LЮ����x����g����	�o1���n9���Y��� ZP���g����Scs(x����"��-&��-�7�u6�����k�h���G�1�ЈH�,��!����s$_}q�}w�Ҕ*?�����^�zD��+J�������@���O���ݲ;�+}(��\�����!~��!���zB�k�Jp�S�o�L���Qd�U���Z�*���=�S��f����L@�W��4�w�_��-�`�����j��Òq�h-�Ǉ�u3,�{Ⱦ�w��r��q����޾I�AO!�M�Jr�%C�D�?���_�-��� ;<�7��%���NH��=]N�����8x���c���ؤ?fXnoq������Qߚ��gU���L5N��7��\����6A'�Qu��x���9�w��F0]��oZ���:Z�̇�U�D
�T�o�(��w[�gp�@��ΰ��9҇
���#���.�'4w�s2e����=2b�-�^S:Y'��/�Jg��7l.�cuɞ�kP
U���s��N[~�:֏�}������1�T�y$�o���_�l[��f�KZ��ze�6�[	~�Sc;R�4h���@�����L�o�R�p��/�`����eHN��;�ݐ�C<w/eCC�ik��Y.�M�6��,�!�Ŋu�J��ٶ؟���G������~H\t*�_Q���ґ��n�R>��!�h�Od�W����^�\��| 9y'N�����F�Zb��U`�i�(�b�Φ�T�������_��my���&|P`�M�P�K�*v善�yź�er��&��9���}`��z�?�!�XhqĶQ�fc ��Лr=<+��U��
����Ϲ��N-�M�+��-�y��/��}�����ѫi���5It7�(' 
г́W�uF��U�q����#�,��L[����e�%���NP�'֖�.���FKԷ�͋2E��O^���z���XI���T���GL΍�&^���yէ/,A�z����ux�eAv�$����{Ƨ���"�~=)ƱE$�/�� ��|�(2&oo�������y~o$[V�%��2�%��A����[DOI�@��8����j�H� !��C�a$Kn-r��-�t`�.Y+�_��� ��������ȘC�;Nv%@!�o(ۯ�11DEE}.��ai���R7oeV���њ��Y�ou���ߵ�v�����Ԇ����o��-����k�5�Z�F��#�����g�[P��{ň5�u��� �v#Ka��L%������њ������r�痊v�	B�.6h
�WK�Q�`�9�-����8�D	6�|���@���_mH�w��Q��2����ƈ����ux��e�E1���K6 A7+7�skq�f�����)o�._^�1ږb�l�4����AK�z�`���0�rn1Q���r��)J=Օ��l=KM��&m��!��b������	$�.I���QXT�1���w�i���V�j��x��B��rR*�'z.��H�9��U@�`lQՐ!8wKWՔ�$cN�+��'�uƨa��ɝ����m�ݚگ�.H@Į}Ք똚�Cgv��C�㱗g[����f���^�1_S�^{]���dw��5W��_��)���#������[��xv��T�-&7VT�Qlz4�]f�vA�J��{Ԯ�G݀];��<q�u3@����!���U����:Me}����C�B�l�����J�!ᛂl����G!*�(�fe#*��{~��U�(�����Ct����� �HH�k��"a�B33�������0��m���ɼ��Cd�gJ:<�kP[n�����.�!e�y���3�!� �}tg�8F����%*��b�����7�zfO�]�cM�>�-���ϩ:-8a���~���CԦn�1�f�*��z������p'?�ۀ�Ҡ���oNѷ2 >�)�zoQ�;�ēT2"J����|���\^b`��Yf��J����7�5:r������*+��+�F�R�t�_a߬0�`��&��|�!1�3���!�,��n����G�o���V���\�{\`hi�k�q�K�!Ѫ����j��:"j3�BT����cv^�.8�H�ǌ������,���$j���[[���������|<r����Cd��ZE�u뽚�`��/���}'�)�a>��s��v�����O���ؖ���U��ꎠ��z����N����b��_���J��"�J�W����m�)�X~��z��a1,��[|Z��-Z~�P�̿9Y��ߪ�Ř���P]�R��������X�3iV���{3���āWk������o�))uW�X��ࠗDd$:꼠��O̬�u=<U׉u�d��Meϛ�&�H��T�2Ƞ� _�ۉ8�MU��*���#�����M�E>��Zܶ����I�5���G����E"�3��c�]��iJ2�o���2?ӟ�\E��ߦ�q1O�x?Auv=�q�U�dUעd�G��\�r��/����M���5i^9^�ݟ��Q�̖ `mq{s��E�o<d��3ݑ����f~H�� �I�����*�sw���9��$�O�x?Ӛ�;�S���pU0�J�q��j����O@rm�$�J�8/m8�����Q�i�|G;#�L���r�� F&����Tw�Ӝ[|����}��lH��
6'k�\�p9ܷ��U� ��O'��c$N��'��Qc=5�(txS%�A�X�E-��`.}Ukn��-���ڪ�)r�~u��C����ׁ�����ؿ�b��x���>-�����KA�����q��.�+�����)��U1��Sm�q)��;�����4;�\��d�a%�Z�O�hꊒ�֗�Lx8(*�qkQ�R�2aΙ�>n��I��ק���*�r��S�����+Vt�b��� ,0�R�s��b��ѱ;3i���+�'�]B���� �F����?�M�W�E!�~������֜�8���,8+=X�P���L����&=M�j�^�
c��I��d�t�[C<w�H��g�僕��[�z�����x����ߋ�����HI���^�v�7To��#\%������SD>�1�5�hee���*w�Cs������?����d:�ު�W%6M��g~��ڢ޹��9�<�8������W�j^\��)8���G+X�����H"��ܶy��B-��rEz�WL�	�,/6��9�R�rM�_��� X�/�^�:n�j����	��7.j:W��w��`~��f��'��[-��������?���������(+4e�8mgV�~GCm~O+�.T�w���a~�%O���G���ˬ�Rߪ�N����3��̇��z����dy��&�k����I��FF��IŜ�)S����)����.ϵQ0����`��f�ă�����?m�}�S�uj"i݋�����؟`"�'D�5�1�$��<:�^�( E����t�d�����b��b�5f��Mt�������t(�P�=X��)���	6�����T�=S�����إ&�
),|lx}�xs�[m�C8����3���C
�Vf��jU�M��[���`�sm��r��b7�*�>�_�EY^���w�7�nj|�Nl{X���N��i!�ǟ�����s��@Q��F�[�f�`�e��b'��L�P',�LS�R#��)�"�����]{V!d� !���_-��+:cF���u���e:��Ԝ�ِB��s��@���'�f�^��J��ճ8?\G��/�/ ޛ���I)�OX������N�����^x�-��G��(��O��@�X�����ß���f-r�o�`�'��<�+����8���W��Y0���u0WT��%��ή8�f�4>WR�������ä,Kه3�ey��F?&��(�JwB�I<g�Ti#_=��Rt�Tx��v$�'�Q��	&��������P]h�����P=��~���?N��I}�X��5̻���J�f�V,r�l�1B��yx,	-$ ��'d��N�$�y�/n���3l�	�M_�M���,�ݼ�B1�W��'����D�.���p���T�C���>���J!�C�v���S��(�Ɍ��7��w�2��u�5&��Z�!?T	���;Bg� A ����[�(?i��Ӣ)����Z����s�:�	h��0�c��~��&���zc�<ztn�C<zi�����c��h*��3�'���/:x���T؅D'�F��Oʹ���E��^E�,N��*=�F��p��k���^�.2�݁�V³(��oS�ܶ���A1!wi����1�=c��x�j�:�C�Z��x�^��������9a=x����A���X��^7���#g
����0=�	�H^Ϲ���ִ�SN�M"�����G3*�Ot�L���E���!�x��������S�z*�A�bl@��a�-gb(Ѭ8�Lp��ޠi#=��B����_Qe�3���#��,.�`TŃCD:�!�|��(��o3K�W�>\}+���K�G��+���_���B�tO�Y[���������B�Z.�p��o�yƂ�M�����WxC��"���xB�49��W�W��<	mEn�����c9=<�u
bQ�����s󌸼�v��n�%�*���E@�����̋�D���co[
pCX,��=�����=#k@'zeWT�!p�� ��܎3//�y1.��&��Yl��m�Q���oi����ʳ���߰�UN�#����bhi>���_�V�f_���Y�U�t]� e�2�9Li��9P@`�A5V�Y7��Q�����O��W��Ab >)�h{�8|^�g����Q6ч��n��f�lY�Y��IIP����d(�fe��P����W1��3/��y��o��rx���apOQF�{�D�ë̇���Do�����N62\���I����g�kS��ëv^�*3n /T[�1��%�D<IUQ�D<�9��!م�Te{�%�CĽ	`�o����hR(}�B�����&�
���0q`b�×�"��ԃ.����#
�?��/�ݨ4.��"o�B�4���^���2�:�Y�1�|խ�6�B�/�lE�˸�┲|�~D���{�Q� �(����lO�ݙZ���Ns�I���یc����*�~N"�z�=�sj\O6�"���=��l�9����T������s�w�o`aV������ �R9cD�a]��)�n��y�L"d�����&_:�8���h�N@{���Yp�f��ч�l��(�Z6��'��3�:�N���(�Zh�K���A�t�j	 �)edḽJ�X�(���16?�&j�
�n����Ҋf�<.������N]~�\�u�##�`q��61J�܈.��I:|VY�-t�!��c&R/$Ȁ�y���:�'-�<������B�XxF��$^���_,]]�?)�W�w� �e|�l�xӃ���}��	�I��Um4�U�LC����߄�H
��S��D�;�u	ݫ����@:g��[KII���� ������`	���ѭ�����_��U1F��J�0@��)狰��|�E�:e	��Df��v�����������E���]�&�e�mMCj����d]�"�.=�mᘘ ����N-1�YHԛ������vG��w��|�SE]os97���z}m����sP(��f����yU��䫲���>7�H��Y,��6K�6����V�����u\Fi韏��4h2F���C_y��gzD�k��K(R6j9@2�/�����}�A���͵�%����g��XIrb$i��{���u�;9�b�����{%�%\�"���1Z�M�ۊ���� 	��� b�XQ\�Q�/��͐�[��j�H��U_<�e*�����+++�\گ��]c��A��!:�������쏄���O����-�E�bh�.4�8�W�>��m��=���'�����c��L]}�|�_�"�<o�/�8��J5���&",�H����:�E��@A�'tP�	Ff�}����+��J O���p�[���4/q���	]7�3aq9��"T�g%��d�9�_���q��R@�چ���^t��ϸ��z���K��i"��l��q���%�8B�yYZ�C0��������B�{���Q�O����bp�(�p=�u ?�Xd b!fIf0=H"׾�aW� ����љ�=v]�PW���ʤ��� ����$}�;,��<�ʕ.���*'	�XL	�T�*���|�T2f�T;�����ڂ:f��Av�N#��s��_@[�M�m��<���*8Pox'�U�4}����O^=���Y�{��}́)�}��Q0�vƓ��4�Io9K������<�"Zm�#kV@
�?y���矼�AT<J}˭wjH5�ҙ�-����ᒬ�8��ae�ǣ�B]�ʓ��R��K��Uy|�����"D6�fsW���g��j����%�?C4V��P�&��ԥ�Q:�O}�@G��}%�K�m��b~x3�nl7���MqG��i��H"H;s�"Jͯ	я��F?�O>l.��<^~28�]���"K��y<2�t�к?\t���Gz��mY�ٚ��R����/+�s� ���n���!1�!�̋�}�5��D��}�o�4Xib�f����)��B��*�� b�$�
2<�3�_�Nt�d5u�e�����3���="��sOW-w�%ۅ�g�s�(�mn�tSw���������x�i�J99iD�����-t�~s�95��I��:\pRs��XK:�w�T��2��6lyJ�vt��K/�
���+�/�����/�|Nb�o|�'wO?d���"�C�=W_Ա�jpt�r��[7��Di�����eaP	ٴ�T�V���2�jD�??�i�LU��Ej����?�����t���Q}�We����%��@ �xcw8	����X�\dJ(J�cs�����h~,-�r���r\�~ɍB�'FK`�gK�A������T�h��`��-'X��(���\�
�n!�)��餪�V�QV0x׭����R(}u+��������o�wR�_TD$���FIw-�0����-�«��W�9p�Y����ӉZ�c� hP�����5ml��T�ת��v��p,��z��l��&djJ���]Ĥ�yMMtCCC��'�o9Ҹ#-Y�8�����3��)�k%�lm�B��n���))5� v~�Wݖ;�0Z��OʉE9}^a��䎚*|�Ӟ���z\Cq�N?�X���Ċ��y�+�Ԓ�hP1)���o}�b���h�m�<�z�Ѽ�F"���O��|�q���&:�m��#��o������]*�ݒdz�O>P��魂Vg�μ�w}�~\j��d���:v�s͕ţ��H�A�*c��?Y	HՁo1�sBx�^���c����M�x�������:�"BBA�x�,L�׭���Y�'�����r5�B�Q����8w�_}�r���́_u���z�mN̥�{D�ſȟi��$=e���I@v!��ܮ��dN&ޢ՜�fȪ'����m�\�
�Tl���nu�?�tY%p�g4��0}~����� �R��[*ܦ�\&w��7a�����e�GO�f�c�48��+�>��?0�Ls�*aـ��u�,��+ޛ6�Y�4���d��7p%���¨~�������	�zKr0M�ރ��]K��CRF)�R�
����?��4�O�o�9������o�n��n ��!�9D�+4��4�)��G#�a:�I���	�r�H"��S|=�@z=��h}cv.R�؇r�0�1��I�k������0��M��*�������������)�M��J�er#����bI�&���#�ϋS����K�b+�{Q#_ԫ��\w9|����w�0�V�d�wުW��@�j]0��7������&��oV�xk�4�u����_�I%h�_"Y��0w���~�m��b!�K��1C��+��e`�3���E����|�	��5��EP�B�ʷ�b�`v�������H"�H2�p�p!>�S���~��z[��X�©ߊ7حd�W]Be���u�7�T#�Xs��X#��
i�Vc%��a�\�X�Vթp������?���Tx־�P�?i� 9��9�'�����/�
����ޥa)�G!,ϒmF�P?���$�,]@�y�+�eQ󡽽/0����-�<�l~��g���57�q�s���={hm�}�`}Iz�q��#4"�K�������T��0��u����/ة�}~&�V��N9qs\��oq~��~D�X�.Ǯ���A�kĒ�*������&�V�;�:#�cTr4���܍���ɧp{/����e�УR�Z��h\����7k|0�ü�A�H+k�z���S��ܦjbX�S�KK�����X}\���|.�T?=M����N��o a��@�7�&''Yi�}O=6�Qf#]>�t0V|,��+�y��>�������18!?��Nӵ���d��n���ɮ����2�Gy1��۝�d�t�m��}���s0+���v�/A��}B�mx��JZV��Jr��$i�W�9�u�,��K\��$�L4���bD�Q�,}�Y���E��;��¬l���Ȓ�I����NLFc2���c~g�B��ɿuuu�0�l�{����_L��͆x;~T.��NON��lc	n�*<����\��v��{�G�[��<Wko�����w�`������Eد<l.:��GjO��J����o5q!�m��;~V�;��/�ޤM��G8��#qv�3�<,KE�ȰC&����?Yu|?D�'#R�����Wq#�c!�� ��f��T�a0�W�0�$�)vf9�:ڕQ��6�� p�+���@�&7�5?O���H#Z��WGe��|���؅�lC�n^__ch3��1b�/�.!PEO�\�l�ͷ5��E+o��tf·�"6��P��|��5���3��}�:Z�>uͱ?�|s�:���|���E���)fg�<��W_�z�L���	��'�,�	Z�sף��.�`߻�#"ʈ��!���0�~.m�9�ß!y�c�^m����~Չ�xO�=Q�Z銨���r:瘍�
`4�ߥ�x��1z�����H�xT�l�V��w�k���ZO!akgf�A_է.՛\��'e�B�9^8��b�l:���U����M]�Bm�p��*����^�
e)�o�ȹo&�~
Wj�g�K�h��[�z����aP��Q�@m_��"͜��I�fi��w��	z��t\ ��#q�y��)��+"�x�V|*@�;��~	>�iY%�[%����ͩ�7�NՏ�k�3��hk�;U�5�%�5dv����N�b�737'���`U�wed�m�>��e�m��rs���ZT�'�v��n����Z�%�M���u����c���u��&�z�,�:6�.a��8�nاD�JL-e�uև���/¹+����̷�r��h�غ���C�j	=�Nt��]�ga�ں�v\�Y���.�骎C�GՂ��3q-����G%lI��S�
Y�4�ۧ;�&%�Ƣ\5�I�.���<З\�ڣ� D���ZO��� FD�iN#�"_5͘_�$u���(����0���\T�G�lX�+�p�/Ow�Yņ��s\��"��|�G�/���Y�"x*����j�>|���Ŏ�@�Ȃq��I� �W�o@�������+�~w�� �i�7�%7�A������"�]ވfM��\�>�3�Ưg����ZIz�J{�Rأ��g|�4�UQ!���Vz�2n0�)WT���������P����/�ƃN"�D*I�!���DX�����m%��eX��Z��� ͻ�ܓ%s�%�u��d�u����|��!��aј5�jF���}�E��H�U��^5���i��UY������%%�L����P������'�x��8�� Ɖ��ts���1}�'T�E���Y|���͌\#��I]ގS ����g����E��-�� [u��ۈVl ��}7NN��1|�'���,�}I4L$j�J�����>mM���ʋ�����B'�T�ah����`�$���_���^o4#/�g׀#�~�A"�n�~,1�2r}"`m��fŒ:|�
Zb9�>_85�+S(���#\��0퍝`�pVT��%�w��
��)H�H�w���ZT����Z�Ԣ�]���sV��yGϠ�������"cX�%�SEf<��ۈ�M���ܟ1���|}�]�B��Ƿ��>��}HKf�@�cNW�o����E�������#�ǆe�΄�*�b���^δ�% a费��:
=ܿ Vd�����(��h��H�qY��nYW�� ���L6��P�I���9q@~bs-!xm���*�e�Ͳ���~z�����7%�ۛ���o?�6��=�o5��2�0���O�>�|�� 2�b��1u���W��w�m~����LC�?���Q)+��r��|���\�f v�$����������>��֍9�6�v2#�?�sv�-�l�ڭ����`�7���|Id3I������z�kGߗ��]��7����G���Y��K8�#ސ� �@Q��y�	S#{p�O^>�!$��r��\<�I �U�������Q� ��T��1�r�̀���f��,,*)�	D��۷yVU^������C�
�� ���������ڹ���2}�c�����V��	y�W��k�&��4���j'�x��ဤ�r�m��">�; �-t.h���c�#G����; �*���Wb��ϊ*�c��?��#��G�u,/`>-H�1O:
�(�9��(E4,~e%�h��z���X��B��l���%�#,��+�Jņ�f���8�� ��ԩVV5��
ִ�V��p���_�2�\Q�ٸ��Q�=�򱺥z+ ����f:�)p�����|�eTUa6Lw�$�i�n�C$�Cww
�ҍ�HHw�R���Cá}��y�o����u����{f�k�����e��u��y�(��<��d�X��Np�[�E��T�d	����?��{����dƮR�q��S�\`@4�|m_��ל����=��6�S�'ϰ<S
-��h�<:2-�%�>��Yu��?Q�������qw�i���q��_ՙ�S1�j�e^���%Ӻѷ�D��9M.�P����}��ul��FX�\�����GGO�V��,̟|�HS�ϡ*�Z�2tL�<��'�}���_�����5T$��E����'��[n���i_�o��9�h��<�k�6�3<��6U�%5O<¨[V��s &�<�`/\
�i�b��� `��J�߆�K��$X����y�fo��7ƿ/���n6Zs4�3�6b���Z�Y�+6�Ǵ\�C겋���umC��0Ye
�镯9t���я�tg���k���|:��]]��JA�t�LYbf��n�����W�㓓h^y_�����BqN7�*7�0ާ7V�X���V��T0{:����a���	�D����dm�wc��%�7�U��їgU�	�
��p^�~<%b��7Kx�x��_'���{��U�)�X3M./��x]��ml��W~�՞�[e'<焾��e�dB|�|�����*1 &x<%$�]	)���|ݴ�AZN���t��)����?Z 5�����묢��8��0�DfX�!���kV	��SQN���A<3��"8��5L5�-1�|�b�^Hw�,e��3�l�c �q9'RNx'�
u���X����{Eϰ�J�a�h����.�ϔc��EVJ?uCGiIJܘ2���3Ѷs�ul���M���%����\�=B~U�� ��@V��B�wM� �P|ن�����&hy??�� e,Ff�.�u�<W�ܦ/OR:bY���xqY��3|�o���5��b��d��'��M�rmP�d��>M&@-Ԑ�I�G�|w����~p�YKpӄO,|g5��TA"A��y|y�!L���k�f<�.�͗y���gz�w�����n����.K
�j�n�9�kf�7r�Q$����C�O��φ<�(�3C!f0�헺L�2��R��}ۓ�o>�0˜d��֗H,�� ,��?!PYE5$�3������js�6�ߔ0v��~<��Ҵ/��r������i�1DU��T�Ř�#�zBB�F�o��gRBn������ƽJ�Ӛ>�'9��Fq�'�ѴC�˼���ׅ*�>�!����O�+2&Î'��<�ܤ(>{���r�V��,�q��"�>��Ņ��`[�D��7!���ϓ֬�F��/)�����l?��g�}N��v�K���]eP]��GP�q�~ܶ�I���M�X�c�6�Rŏ�(����Ē�����)q'�Ii��X��ؓh	��D��W���~�F{w���W2?䙂vĻ���z�Z�������V0�!��C��*�u���J����za3��}�����N\��&'�����*|6)��<i�V�2�"�bA�&�?8�� �BW���~lm�+�\6��o2��V���1�<����/�o~繯��|�+��,����R��g���h�	L�\7����8�s�?o7���|��� �+�`��JZ����.�Cm>��/���kI>�n�߳�7�������Dp4�/�^h٠�� .Aclhjv*u�K0N(A?�5��2�u����Ӝ��J�zfJ�vhZ���f�iZ��nyC}z�����^��Pf-�w����1���m��b0j�K��������t���v��{ގe��w�	7��4Ьȼ
߆�OOs����	���n���M5�@�=?3Y�ӭ�&������kc 8<r��*�(:����Bvp��*�
7��혉�4����ަ!oX�is�Q�\�ا���n� t.��Ǟ.����z2�u�V{�Q���X�i����M��=�����,GD����d��PB�f��s'/��v�crjj��l�P{��������w�U����2��NF�1��Y)L_t?�69[ȕ;�`aDQ��:��G�^�����S��U�ݣ�*��P��dY��G>9��}�����>X/O�����͛����Tv� =�7�}o$]廃���W�B��w7��Y��> �|�n ��f�{
���v���������8aݞ������z=��0���b[�\�W}�1��b��L���_�߳k����QҐ��n����sb���X� Ot�^59����#]�T���߮�k'�|.[�uF���]u|����Ng�����Q�̕�},Ƥ��>&�������e�#�>�E�3*�^�-.|����/��6h�������OK�_���K�':�8���p�nڨ����Q�z�(�h)����!g�$+1ƷL�o�5�rot/ ��'[-�S���2Ja��y�<���XW�V���^�x��҇��q$�d� �=j4�|��-��|h=����c�����kjhl;d����CS��g"��D�_�/G�4=���j/�X0�(G^r��]5<l��~I�#�P�ipEiL�����'Q����/
2LM�����%_��C��OG�4����+��B����TM����P����_�p�a��!5�>�N�W�⿖��4@�.�󫈛j����Sm��?N�GQ._~�kyĲ�����p9Sd��N��?�U>]g��	E�(��dJ6$,��ǫ���/�m	#*Ar2����r%^����B���Ɍ>U�>)�Nr��� p�L�N�{��lrɖ*�����2 @
��d�F�qu����'{(���Y{ZW[�rL zr���b��t����:�D�"����t/л ,s`�6�#&�+=
φ��D�'ïuy){��0}��, ��WP��@��?wn9y�?�#8���/4� $M���{�/歎���eH����?�)��7x�޽�o���g�	O���z���+��S���䁐q
D݇wE�0x��NBp�!E�Y�O�c�N}:�E1�g�$��m�1͸5�
ޤ�Y���7.��Wl��&����W���D����������z�5	�c�m��1g�c}zi~>�~��t���ѕ/��{���Vo�D�K+����',z}�v?o��,bwdќ�N�Y=x4ǮI�le�4�5�~�����C��֏���11����;�s~����"��|n��J�� ed%�Sâ$/yO9n=y~ZF�X\I�齗k+�4-2!W$�´�A�V�G*~5�,cY��ݙ���{�*ġX�~�+�����G��3D\�P3�����/�$_'��#"8��q��� �i��ܰ� �1</@�VMc��~T��g��jy����'���g;Pa���Y��%�Z >30<��i5�����!kK���MUt�<�
�]������9�h��}
נW�8��qҖＫr�:�#5�Xb����pV�U?5i�ʔ,��e��c�y?�����}�ȉz�רZ�'�2ؒ��?S�
�BZ��w��q�߮�-U�(F�+aӶ�E��5&�����|��l~�M�Ǫ�vz�<ն���&��3>��
"��������D��p�a,v����iA|999p=_�/�B�,��- Ɏz����k����O\�ݧ��(����&�t�C5�A��%9fb\ae�d�������-�R���r���ѥ<:O�V�u��N�z"��}�	�*��bλQ:�.�����`ko����u> �s��u[�[�׏l��wg�MM�x��O{���YV���ވ��SfYw�P.�
�v�w�)њ-�ּ�z� �X9f"�:� Gc6��N�T��Z�-S��b_֠Aj;v��h�?�bH�B)D�`f�u�p���M���PT�D:DM1�7>(�z@��kX9�76�wjD?o������ԧkP�HxJZ�zݫ�%|w��g(S��O������x�}
4��#,|��@�`F��h�YW6"����Q:_�ji�!�ó54��l��;[�e5�j]<...��#S<<<�}�"9b�.f�]�#D�������1����(�O���OY������ƯS��7麸�u�6��#������S��)���F���Q�Ϟ��U����&�L;�̼u�/:^㼱y���jX7 ��,�X}�m�}����$�;��jm�X�s�8�����ln��'nSv^V@����vӧ��l��;Z�B+%���R��z���rX��C�����7��%���,��x�>Z�Y����A�bWۗ���2j]������k��rzw'�޸������x�\=�d˧F�3�s[t�tg�q���9n�,q����D��:�����M�l�_W�#�:��<��ӴD霹P��`2�u||iyYE�n�sI��Q2����H�+���:�nc{P��~RB0�w�<2=;?��?�U@'��s�m ��'ͦ���XQB �MTj�y���<;�s=��k���Ч��sP���v��%/���)�.ki��-��>��r��WZx��
Q0N�����=��J���zF��hԞ�|��ۭ����^@�6����O��a.��Ŭ��c1���{0;u�e�,���5����$���	��䋋�T;��n�]&-�*	�L�����ځ-�j\Ѫu�*�� @^��_�:��P�����I�xv�>Z���Ug2�l�f����/��Vu2�[8)�ql5����8XX��s?֤Bcj9կ�6s߆e��|�_��;������[�BH�Ȅ���!���e;�~��O&ޚ�;Y��c�����/?��퀯���{���Ѹ"����t@@�¿l�~ߙ�����i�P�ceXJ��$>K� �,~v�T������\�Nt5�m,�0��f���q"z,��X�K��J�y@���`��!�J����Aw���6��tt��,�j�Ƈ�ŋ�r�[i���zE�EnRw��P�D��=�����!_I�d"��T���""�<#��WBN��=Q�eN��X���YX̴7�}�@�*li��FQ�#��7Z�o���#��W�-�u,�S����D
�<�g�no��`�.�2�5���{R�T�V�~��9 �Pf��3B�L�}zz��qjq��p�>auJ�=����w8^�6�!�+8o���K��(Q��ag}R��hk���c�`Ϟ`�^�� ��Q>$0�*�>���:1AQ�W�q}}�x2�/>6��������8yT��୭���,<||��Ck2zUY�[��<U,F�q	�導��Ƴ��lܰ�.���RX��Y��<��`y*�RV���%��}"�D�׺�|��R�b���qcXl�-���k�w�bqryMMT@�;�,4�9QX��D��/��}��t�@m���˼O��s���&TP.oL)�a�C�;��h,�~�6�Fu
���&�.�/�O)�����؍��$�D_��cK�`���4S+0��y��Uf��Q���h�l���$�҅rĽ��uR�w���|B���lu�;�^.{@�p;�:E�?���i��V�ߌx�U�1������I��1�j�!�)�]�3���YP���#I�j��eNV��7�#�h��Ԏ�|���5��h�t����$�(a�u��Ky����`_SK�ʊMTL��r������p��r��lи,�_����F����YX|��87UU��Xk�gՌ����Ja�f��|���סMKy�������aT<�V�T�L�̞2ΏB�?���[���{�%�w��S`"*7��Y<��J� ��ayy����6y��/�)�ttt������:M�A/H}��G�T�����aU�x�*!C��X����
~-��pՄ�V�20d+�@O�Q\�M���C=�A��D�&�H(�&r Q�˽C�|��NH��7Yx�I�F�D��k�v��ז4���IDŭP}ʲ7x���`w7;��K��S��H"��|x#���N����$p[�o������b]�"N[Q?���Ґa�z����"���Taʜ!H.�[~�6Z��P�c�>5��m��E�Vu�5r�8����C���9o�����t�p���,���Z�>|�Lk���T+N������ؾ{SW � W�Sq��7�`[���6��r����N#n�ԱAඬ�`��.V��ÚĮ��>��g ڃ2~��f�U��lB�iM~�(<~`�#���<Ԡ��+A�C�
�2~�st���f,r�a�=gDi||m�f�;(Ң;F�f�=�~�K�9|5ۼ�Fb��Q�(������3K*�X��&���[�%˟g���U��#�-Ǜ���.w�R[�W�H座&��===��n����Z���Q���;t|��Xi�9��/�䲍�h���~���w���>%e�:8�ޤ��"a���S�
�u��5���WGK{gUXD��%��/�=z�M	i9Vҙ���P	ƻ�\A�搰n�k�>3k�rhXߤ���������;�V�*	F�����<���iI�䪢"�Uf�[OmV�1��k+%��Ye8��ȅ,������g�T�Uϝ��\�ŕ���f�:-(�s��(y�jN|������O�UΛ�b�4E�RE��em���0�VnK��ػ�s��=��S�ӛp'A���Qt�㭨��jِĘ�����;��_F�j,���C��{���;����N��^���^��
|�w��x���V0b��A=Ekձ%c�L�b��`�%318�����@m����i�B�%{�ZZ'ڠ�����̟��6o�����UNN�%s�J�[Z2��.-UӚǡx�P,�.�}��_��S��wA�pX6N䠡 ��$�V�;����q#f�%��n}C����.��ض��u���g���w��bi�jo3 �c����I��("�/@��s������6�^ŭ��8�"/eo�g6>Aa�7 ��ir ۃJ@� �d��_2J^_��]\h��v5���9}�	�{+D8y0��v��+k��YO�8@׾�ӾJ4	�u�&�I1~{����-��s ��y�U��C��\��@�T�J����3Ȏ����^��yE���L ��lP;�8���{�i��18��Ih��\�_y����DC��`c�7��<�����[��@G�򖊜2= vZ�N{�4���E#>�O�#�va	�ܜ��]�Ki�=+c�/����w���ވ��G�'�7[��
�{C���t�/��E\@>Ń&{yw/��j|�W�xL���ϴ�e���ǨY�P[;����Q�Lu8��A�C��/�Z�E��y.�,]��ea����Y�2n���Z��хU��/�Cn+���'��8e��m�A��3�F����IB����y�6�x3`� �;8SHw#���Y��Ǌ��� ��ʢ��<b$�At��2�K�!� ��D��OȥNt aNP?_~��qj;���d���Ťn�V�ex�A�Ņm��S�����j�s[��橚�� � ��n��=Vs�ws��Ǚ���$Z�K\^�[w����R�K5w����˼;a�vc�3zS�8�룺r�wZ]Q�A	�	���Os�L����U�q5�3i�h5��Ldx����G�ֺN.5���+�����ݠ  Z�Ƕ�ܷ@��SaS��ٸ���O_5��x�@�(s̻z������43�Z9J���+y�u�rBڻv>�/8�VDx�Iz僜�i0�r4��l_�c��0���WTV6�u}�H�R̪�wĿ���9<�����W����,�`$��'RI���1}p[h�UǙD�lg52U�JdMud98�t�	}�DQť�����ag�6Y'�+���P��d=��\��&����w�jp�=8��ź*?`���:v������t~go3=������=#��4>�mI-g��ӓ������>"·Ԇb�X>]��z�O[ ��!�M�f�"�����'��KX�I��u%U�'?=������V�t����d�
��ހ�a�~�����(���\`��l����IC
m./��ס��3>>��}�~����x�?5�.��S��8߉��8D�J�]�[��0"����/j�P�֟�돊����W���Z�TXi��Hs�w´�N�_����;u	�	��LLL�������
a�AT�/??�*���B��
�w������_D)2[��]Bf��>h3�ե�r�Ԣ�E����V���um�Qψ�vS��U]��i�KC�y&�5�� qͫ��" '�q{��@��o?+�Y	����8����#�'٦�ǲ�4�ػ����^/����.����3l|1��@�!�~����n޲�� R$�f���?c�}R��5�;�Yis�8e�݄M--� X�ˠ����6�>6��5�P�?r���S�<����d��p���N��H�U�Wc+[{b�2��߯�(M�^�Ri:��3KL��R^4�H͒���(�~�9B�aI(p�����wz�!w����4������ [!s��m�_$5M��Ѭ � }��QIĞ(|����g� ��|�p3yp��w������Ҭ�,#�E�dZo3A�ë'��e�֭�������lX姹d*�b�/�ܧ%ˁ=z�����;"I,b���*�����P�{�!��8��b���@���ǲ��w-��6%']�b�(#b�=�V���C0�����w�o6~kѭl��O���k����v��WVj����bU��Ѓ���q&� M�Ծq,,e���.�'��$+��6��CT\�¤�V��l�
m����Րq~[��6%�X~�I���d�/�hx�"�Z�t��{�y�2I����@Mw��J6A��'�����j��Z��p�)��)"��KF�[���;R$���X���ς��*U �&2���8�{��C�ZZ2RY��/߼���9=}lf2�)�r��tn���=G?�^�G������א�8K�2}�Zf��ld���X����"�2������S��wD��ˇ���T��k8�3�����cV�(����y{<p��s8Kj'E�p�e��G���7ԒW�TQ������<!b;���Ō�˩w8J���xv�g�Ծ}���?_L��;��Z��8I�;�bxz�ȥ���I	��	�(���k�)>^X
��6?������蜌jS�Z@��U��@3�!iN8$*��o��-+��\{�p�c�V���y��ț�6c�w�qO�^M��%���r� 1D�J��&3���^��i%<�:~,���"�.M�>�A䲬�|
�>~ȏh���7и3��jҼ�Q��|ںrm�!X�Tӹ�[qY���!�߽�� ��n!m�� ��ht>�'%�F�L������	�����:F������WxŪ*�N�+��D�e��VNn��WD?��M��ʪ��J,�W8v�=��ܓ�2��u��]��>`���6"F�&��l�=�xd�A3.���˚Q\$xd�
F��8x�__���}%L���H����Y�2�f�tq��J��GO(�/��L�$/'��ʞ��z{��v���z2=��wY0��)m�)�P�X����D
��.��?+�b$��~��������p���������K�ȭ��b��#�kh��[w3Z~��-i�-��V��{G&�4C�۱J���j{�*�NE��j_��2�t�V�XT����_���|n4��۞ڼ���Ӆ�w���@
T%e�@8��]��*(�Z��e�yYM��)`��I�r�8����Z��JX%�9���DGl�y짬��[������ʹ}���H-�m����ɷis��{܋�}�U%���}d@e�9��۱��XZ1��2�;���0�og�ķ2E"F��Ix}-�T����F���޳`3�B�֓WM�(�~������m�5}'����_�߱wO0qʓa5�	�nps��枞ׯ^�yq	{�X�|~	�U���J�h��V�f[���sa���w��y����]/���Oe���P3^(n�Ɍ��/�6�`�u����&X��g���)	���`�'�!����v��IMg�$����	�5����O-l�R��U��1��f>�Q�w������V��f���`)���`�&�����v�#�q
����Y1��,z}W�I�.�m�Ky���?l���*2 V�֣Lx#s���@��~5�v�W)DFG�GH��H�_y��L��ޟ�kq�=��p��[[Г��>Z	>�;<`��d��"e��|V,�y�B!Xې!�Q���>l�}ơ����,�l�uܟW��2��� �"��E&ZSb�/�o��V�9}%�Q���S�����Lq�����t�@��1/L�:D,� eߵ��|���YZ��f���|�_��9�����;7���zn�~5jN�0_'�b
5K����i����T{�0b�o��v��@�*TB�,�1��2:��=��hɯ_�x��5��(I��zg	�?�ZS��l�4�j��Z�ɗ��[����d�1�8)f���7��?�R�r>��=ف��3)���������\��W��`���Ad������w��/��w]�/:���għݼu�B{��w6c��Hr���>�*����}��$s�ٗ"��{ϣ�4��@��lFF(�k�Y�D��u�s�\v��fZBl�Sm�wpA=Ϸ���l�g�hOо!��Q������)�����I���*H�������D�i��]�!�хO心��F��p
i�� a�D�W,B����P����2��Q���R��Q�~d~{�e�R�Я�'�ML1���-��z����؝4E�D���(T@J�<v��<f��#��{�kr�mK�e���&��%�4�w�%�"���	�F��M"r�T�gxʸ�?|ѣ�3���Z9���a��.�b�U\��������~J.� 9*g�y��q6��K����U��2��&�G���9biho�����?%���!^Aˇ����^����lu�4�YO`�����O��
x��������ۮ�:󛗟�2�ajR9�ͳ���%�
��SL�������Ir��k"Yc��\���`6~����κ�U	�,4�ʆ�c���s����d_���M��|�����X��/�J���բD�y�7���۸ﴩ���أ�Lux��������x�2��l�j{^������(<��R�@M{�a�QR�/z����l~�|�6�����>D�	Nb@JO��r�ui����S��Ə�P������<�&��oL0���I0}���>{�U���K��31�_@�3ʓ�v��-I�%�#6+���&�U��j���a��/��\�*���J����m��\t��T&��㏱pL�vrc;�Y;���#�c�2Sm���o ض�K�����a���"v`=�=p�7���� 8+~~�z=��V�А�a63P�yM�sq(��ny�Z�����=;i��[�?�����Q���h3����q���Y���y��$l�֔��_��L�.�D��M� 15�ڽ���bd�ǿI(�^�#�����\u�e]9xr�0j�3��LG�Qb^�
ݤ�dt�ʞ=(������&O@�==�߳�`e��?u�mߛ��~�iCL�}A݆!��҂�Q��	*$êߵ_LX��4��6r���Ծj�����H��o
�խ��6! �*#� �N�5%WM ��	�
���_w�/ہ���f.'G��|ZBhj���������P��x����{�ygۤY��{�G��he��Pr�^�	AKK�q/�*x��I��^++㶟f���H�;�Z��f笭���_���Q6�����3D�'�8�KR��X�4ʛy�CNi�wEE	�(�x��>ʅW�����t� ]q�]�JR�ۺ�"��qk���-���f�<�dg�j���?����4˗�R�n�?UA}{W�p����(��o�����?��F|+`DRs~�o�X���;=��k��+�?M|a�DGVf$^�\�`�=��0,�%l wQ��b���Qr��-[h,�!�����������-I9@~�­<'��\��xț��ar������"��G`[�W~)GzFF�� �/��qO�^L���_bk��&�
�������H�Fx_��]�i��9	��}ۯ9�c�c�pK��@={�8��K����~��v��qƼ�ֺ�Ož���-|Q�a��~qʭ�6������df~�A��^��mR�rQOՙs���'��x�<�!�f��ID��<]ӯ����tB��nq��Ч88��i���S��$ �2SR(Q�6s�p��u� ���Đ���S����yp;hI��ܩ!��X�U\p�ξb��og����c��l����1�J�8���W�Y�@�Λ������/ځ�Y�b���VdBz��h�,�HX
�B�/����QY��+�=��t�K��tUܟ��&^i�ݣ�j�.{�T��b7�	�}����O���N-,v�z^��u���u6���:z�ôs�����A&�ǆw�%�YIqV��=.0���(�� g��|�����a��foCO
=X2C�5ɚ�2�YP����(�Vh�/��$���!�!G+�1@(C���9oX�n��:ID)Iæ���X�D=�m|\�����s0�2|Z�� w���J�p�a����� �(:..._�k���̓�j�]e���W��Nt�t�p�P��?�����Bi�S^�0�Fr�d�y<p���a���Zn�X�*,J�����ʕ�T��?�O���y��1��+Iw�j�ņ���?��>�եd����WUou|�ۓ?��p����)�!�l��1N��o�\��)1�m�M=�±���ò�4�����Gp�\�@a
�i-��|���PxӨ�c˴x�O���-�-�7�^=5%~.���	/�QW�M}���	i	�����ZD�缆
-e%�C�m2C�ƺ���6]
�<_�J��ň��oU��@�b ����ye�G#/����mP���E:bø��L��S�x�1�e��is2A�s�U���C�@	j�vɺ�xu ��1T�E�E�5�����$����$(5A�؅����������������p5M����,ȏ۪^8��h:q�:Y��&� ����b*�{��Sw��xCju�xC� 8�N�=����SO��������1p�S���,��G��6~J��V�k>m���&9���ZTbF�2�2�V%miQ䖼����Z	}�x4i-�����I���8W�3�&���U��z$Qh�7�����TY��n�Q�"��<��Yl�A��G��M�l��_m
o~� ��&������<�4�����	U[]�G�_$g|E\���EܚF����*6c#%�)o~��f��a���l�7Aԋ҆������r������̗�@�=�Ç>qj�+I���M1YK���W#ÉG��
��m�&k,�9n�9����5��v��X��"R^hԷ�v|y)���:�>+�R����A��=��������y���z���J�y.�����0Q~$�s�����>L�F/`�!���l�E2���ѺJ�JEӌ�Cǩe�����D��$8:�����͘]Kz0~�)��Ŭ��?�����u=��CW2�ه��G7���Gϰ6�/�o>��]��j��%��j5��F�M����]�.��$�u֠��c�����K����j�7�2#'٢���LIK?��g���.��@�ՒZ���c�5�G�HV�J't��ilF4i��� �5�����S^B'�D��/Bìv����'� ,���m&��m�C7�9mgy�X �S�Qh�p|���v���쬫G-���X5Ҝ�5G���$��2���D�l����}���)$�Ȳ�Y�\;�(�p:��(�I�zx�;d���<N>ȋ�j\}�_<}�z����kQl�8e{eu���!��5�$�׻E�9A�D�����j�^λ$��O-�t�܅<x��˜y�~���R��[\c#��abܧ���+42���J��/$��f��<P4�e���\�8ON?j��S�3*����5׳���z�˲�kNpCQCC�Wlu�@�/Er�U�p�l�lAf��SEd�o��f�q}<����H&ِ�Y�6��~i����mg����	-:_w})I���dH1i|].>'��h�L~<�x�J��� ��UBv�.���z�1J��q��]t4N��q����v��'�q�ol<�Ȕ�@�v����^s�<Ӫ�KM��-��2@t���[8/n���H`鄑8j%�З����(��]��P̖d��ِ$1��U3[M�"���<�R�"Dr��}��I�u��]:���\1��%���1���sP�Z���� -ʘ�Hw_̼�tZ��|�Wj57� ������ ��M5%�BP��s�M+��&΀�)����V�S���=��a�R�{`i)�ŝ��-:^O'�u��?�[WGfhh�4(�ؘ�4�ǣ1��{�e��W�Ѵ�&c�Ke�i�D��'���Wa?��_�(`9IczȾ�V��1)�L\�B!���*snQ��>h��a�]cJRkE�Pي�D?�˦�ٙ�VQ��>=L��7�W[���9���!6Wz���'�Z�wM(�j�7s�MٕRY0��6|:9p�Y|��O%?n���Jg���i>��<���zB/Y��J%�,�缁;r�9�y%[=;��~���῍:��5���I�|����A@��p�����AnP�<�R5(���͓�G��.\S�y�H�f@�����L9I��8;94�$��ˁ�Vz|y��r������v�	��=�L?�cυ� �Fi˨���^x34j^@�o��!�G�j�	E��Ȣ,��*VV�N��z���q9'�(DL*��v'X�CJ�T��G��SW���Ō���U���+6Y����[7K��>���k�iT� S��t{9\�����^�r��r�0"Q�!����ͧ�$l.��3�E��k���	/t�2��"���a���d�`z����mL��(�{gW��~�l$����>Zխs�U,���(�5MQ��g��wy�q�E)������F��Mt��U��|����I\پE
�	L����N�zB�{��n������C�c�M.;����/S;;<p��1)|6<��%:py48F961�FL�~]8j3��փqW˪`�|NTggKv�T�2^=�8=����������Z���i%$�c���G��v=�zihq	;�k� hs��ݚWE�S��5����\?>v�q�҆�����J�*��(�"��������C��3u���|���!�/)�5�q	��[��VJwf�s1�1�,��d~��Y
پI`��2�_M�Z7���!7m��V;��%�F�m/�G�0{����L[��@���{��;ѕ�3��̵+7����vA'8��'ײ��>����4�� }V�RC"gjH%~��[c!�nX�xρ���q��B�3�n����̺�ϐ
��;�n�i�1�E\�����I�ͧ֑��@l��^��	����L�I��88�[V��l�r�]�BZ�.�*C�h��gK�6Yn��,:���O��=���l��\<F5�)�=�g� s�����3:8}6O=���N��?&՗�����*,Ϳ�lӪ&��I�Ƽ!��|ꑒ�W���I�*J94OS���.d�R�5m��{Lo�;�h��X�,#)M*i�i��F�頛A�F������Xl},ON��l⭁��Ėo�z�a,0�1��/m\�����<]��6i���.���}��d��.F�&팸:�\���*	J<�-��7��D}�R���$)�A6�FM���u%����Ew��.��+��eO�:�&�V�OjQ���=O~���9n�Y1A�x�R��/2�l���ُJ�Fڝ���$Ɲ�;��;�g���A!���q.
E=�A\Ҕ��(�mp������٘�m嚻���4�_ȥf�/F�jx+�����\�졿�nа�����6���C�#�<���v�ZX��ɯ���U���l����D#�g����i`I[f^ףl�=%�Ɍ2a�_k%�ӫc��ݬ�mY܅'=����߼T)ר�0���9�yg�����%/9����%d��*���7�no��/jrVA}4������V�e;lHu�����1L%z���$��E%ߝ,5�bU��[�T ����c�~%���-c�c=Q"��8):��ğ?u3��AA�f���⦿Y��9��Z�Nt��5�|��8/��
CJJJ�'�7$Ǯ��E?��ywV0�e1I;+�I	��V�^����{�5<���Qy���a�=�Fd/��o��Vv���|�1��xo𔺯P��Q���L����y+D]^��-��^��S���V��k�:̅��ւ���l�`{k�h"�T��@> @�UP�XW����G{:���#�3WG�Y���{p8O��K��?�+�W�R5̻��;�X��-�X��_���Z�i*���ݝ����jqn%���	('.��M��2���FC��FÐ�u.���rt9��ye"W�:p�
�UP��~w��Ck����VB
_Ϧ߅�
?�B�m�eQ�0R4���r�,_���@2��S����}G5\לM�1>F����6����X��6ʁ��V�w'�M���z_�n���i7������n���Sb�����n�Ut�jX��1F;���b�����|��n��]�s���&�)U��piƬ�����YB����k~�����<υ"�L�����ԇc:�}#-�d6ߴ����fv�h���ܹ�Ff�P�HǑy�v=��S���h[��3uR*-�����i�J��5r�J�}D'�	���d/u/�j����(��v���3dد�ã��˓�[�*u'^���2,���A@J����	����$��n��e���A������������.x�㬵�>k��z~��yI	��C�iD�RY$�bu��ܜ/"�/����Z��e�o�қ�lM>l^i�,�ޫI>�ն�+�ǭ�����������6�j��o<=?����\���dp^��쑖Ο��]]�0���T�z"D���|pP�����5�^��{w㔜�6�@��8_T��
�����=<��p�f/����u��;�U�Cv�l��\3:cxؘ&�B�;��͑��������na9ws�qG���J��bٛ�e��n�0/�(�dqG��H�`iǐK�n�����p��Y�I�L�XV�2�}�0x�Nm<�.rx�O;G��;�j�!"!�k+�~݂�0��xU"Y�E3�kx��81���ȃɹ,"
m톶B�1���C��s]�j�|,dh([��<�:�7QV�CQ�k��+g�$O'�.*jy�]�1�t�1	�_x��߇p��y5�[�Հ{G��z���|7�oC���!�4����C�H,�a�kļ�V��3[*��J��~��3a&�����7s3��
w���җf[�!��YL��kD����ܛW����i)�!0�r��is\pMNE���gjP�ýV�7�}�U�|�]��j��&�m�˰`��u�X�ڱ�G>Rz+�Fc'8ϊ�:s+ۛ<�8p�9A��ڛ(���Af��畾CeY�zw� 0F^�4|�N�{�y�T*qlr�%{�V�q)�:�(=����yzg�F�G��kJ�P��K�>�v�4Xd��e`}6X�Ou�7��g���7�VĄ�����&=�7�����K����<!�'5�a��¤���o ,]�����C���3s#���7�{i*���� b���[b���o���hW��PZ��_G\#&�̺��_�/���mh�6�k�}�	�7g���`x!Т2�Hj��!��൤��m��+^O ��E��$�y@@@���F��y�ݟ�rQ>�hiko��Nԉ"��<�����R������0[�;0t:�����ygR�,��W)J�rka�?�lq���+��������T��"9����o���xB��j�sG����ׇWs��U�4���HJ&��E���:�E����w3�#�c�YK-d9j1�S|��[g�J�w�֏�t��!S&�.H{5�'(�"�r=��D���!��4po���͇�=�]�q��13�aA\��.�;�����>�'�e�k뙧�� ��uE['���7
B�X�"Ja�3�1b�pfWB�p��p����Aw��rS�k"�˽�$��r��;^�Bu�2��h��f�D��ui��~��C�B�YI�i��@
# /Evx��Z߰WlӪ��=X&|���d |4���9�$U���W�Zi�����I��y|� ����pv��,�0h8�n�.��n<d)ȿ�����yJ@J�)Db��lw����o{˪tX�8\|��C������4A\c�����Dm%H�Û��%�y�*�<ǌ�<*`�K&�~��y���L���Q���j�����|*iG�<��H��E"%8�����C���	�	��G[y�V��C�����,P����4�O#~C^�(�7��h�q���Z���a�I�)�(������c����ɼ�ɨ��-�W��pW����ڊ�_g��2r���|�� �*[�����7f�c��Y2��e����If�c���T�-�;
ƛf{2���/��2�-���yuY<,�Y՘�1B�3,��y+`�	�e������;/�xx�N3ws���h��B�,i��c�\�;;�&! ᇱ{�GS����[�j|u�Gǚk�};�ܦ�<O�
�F���=vRh�)��M��ᱚX�kҟc��PжR�CKn�2θ/�Q@#}n��23�[�G���A��68��b��L_����Ӫ��d-5�A�2�	�Tϵ߿��ՖK>V~LđQJ����<9�*{�^��|_]UQQ�%�� �0���Y��'{)������Op:�����<�����ú��y±��)�W;��Î_#Tn�:Z��t�
Uh�I��"+������j��$LZ���\j��� ����	��?Ə�9�kMn_�P�+k�^<�r,M�]�_@PoB��qR�DA�b<�`*Lb&|?00�<H�^?H����k���h�:\9�k�e�����z����p���M�Q�����v�ͥ����Oz�K�ٺ��m�׆o� c�$�AdS'��qӰ�&��X:,�o�A�IfM�F�-������%�,�S�!�`����0T�T�Y��D(���'�!��S��ي�)y+�gA��ݖ����hH!�ċ����Ra��h����$P�?C~���Z	DX)w" %��N�*��H<3n�A��11nƑ��k9��[P0��$Μ����#I�]vHcӳ��a�����X���E���<����9 K�U��I���r!ޔH��n�4�+S@��7^?�q� �6L����3��p��ǌ�q��aG���F=a�r߲��2]ei�ql�1s�	����v�>��"���s#� � �,�YYs���������dU"�Wo[���WRq�L%$n�6��xt2��$%#no�`N�yq�!<�Z&z�6A,���jc���
�%��+crAf��V'�͢^j<�e=��_���P�Ǵ�B:���d���?��o"1�/q��q��ҹb��kJ���{$V��ͫ(z����'O�J�M�[��*'4Ī�� ��� Q�BlT�i�5���Ս4C���+��a�>�k�"���S�P��ZւQ�j���Q��y{"�����w	�B���n������SOS�(SJXE?��iy3r3���3�a8���?NQ(�ԝ(�YW���������"x㹡�Y��G;[�F�y�~$Q�4�5[<��^����'�������ٽ��S���x�S�����K}���X�����܁�N�;\��:��a�#����<-M��,�E�^���^��Z0T�����= ��ZZ�����֘rYE�cȨ����&������@4����������;� �p]���oL�6�8�q4�414"��\y�<6k��yjzm���Jy�~6��C[��B��~�8����ʸ���{�:o$�1~��k���®�D2�����!jV)��Z;�KNX��Vȼ��x+��V�)���� ���,� >���뵄�����(!�� |��u���%��?����^��¸�6��P �ڋ)4Ԭ������)zªG>JL�SR{\{V�2+�~,)9�65��{��W �lEUU��"Τ�椮wt���H���Ep�cZ����z���f�o�+�O�9�\+�ΎEI}�>O�'�e*�ij��Q�P��Km�� KZf'5�ہ�'���π�/z]-�4R`	m��뛟e�b>�'��a��|$�u{�X/m��,A>�z>���f�<ޟ|���{;tN� 	����Jf�ۤ��UV�,�窫���<� �NkV��I �5�E��,Ņ����x*YR�2`vG�����me��k���0��~ٛ����-�S�f7K:5o��[�:��>8���p#K��\���~k�L��\w�1��
�����4��$�|q��D�S��2���m�o�TaNE%k��]�eҀc+�o/*�]#sSѣ��tF�WO��<�&��b�>�av}���<��R��E�T����q4b�;<P�ԉY���97K]p�e�o�_s-T�c	�}��%��b��8����,j����z\�?<�?�����y ���sv�"�b���;�8���;5Z���a�w*�f0���"#/��8
�A�'�
	�{���4
�������-:��I���d�(��M�]�ɦ]h�Q��-S8~u�(���ʓ��Y[����Z�L�"o���I��w���ʾ.`ބ_c�>Q���L6��!�c�B��+��3Ǳe�d��w�4��Z�Z?'�3[�Ωab�j�zQ˄��d����>�gK�43ߥ�~n����d��OLrk�(��ȫ��I��ׇ�?�"������y��x	�;��۵tXt���f���$<�D$|��s(�f����v�roez���)z���Sv^�败�ʗpv��=���+�%��ǭ�h�KLu��c������� Gw���YB��|*
��N�ҍ������q˻�S�M��n�dٜ;0�P���;�:o��9��<��*�Zy�:<��?�1����H�Y����mM'w�����2R�D{�u#����\������B��n�w)�zY�/bu�3_�Uy79'�{ﶪ���Rc���������[Φ8rb�$���'W�~����P��q.*R�����c�ڳ�G����Z��2h#Y�����=��T+�Õ(=a��kzrA#	\�@!�z�[|�^�60��~��a�f�"hL��R��o�����>VTT(f�	�J�m�B��yr�/�\w���i���G c��nC׈���ν�M���B{��X��ޯM}j\2S����ٿ��_�kcd�:��g��ml���S����T���qS*G�v*Q�j���]�q��uY�;u A? �O6kDA�j��ﾉ�d���q�A7�<�ڜ�Ja�����V�i�Y�Z�:�]��+�S:��Ӊ5U��S�B��q[l�Ta~���B�S��_�n����|��5cK����j ���f/  �5���3ı��;W��ؘF攽��_������YX�d��"�˸.g^��n����ŋ�{����{F����xi|�Ъ��m79ظbXo��V#W�����1^�=x�ΰ�N���O?uu�C �2&-��1�i�c�c��Ăoo7����!UUU�Qr~-�_)9����s|�"zᣅ�
f~g1&r\D��_��ߥ�w���GC�'02�iǽ�^��K�ra��Ҏ7+q"W}�m*�@D_DF`_�S �si�J��R%���Ɖ}�,��e��u�n^�G/�åN��d7Oם	r4�tq�}�j�M��­�0��-�I�����7lQ5�u���D��lGD��2�p_�0r�Kԯ�+��f�Q�e9�v�-œ	m�6��B�����/��q����ty�\d�Qo���D�r���s�$��ڔ��@���6	~������Oh�Wh4�(��0С��}'31L�깋�����[3�,ֽ׷�O��Sb��
�m-��B���O�||����g�2tL0b&j������f:ݲ�۲�o������o�"G?
ƅ_T� �_^!�P�h���S���>������ήO�Ϩܡ!.\�2|�+��(�����46�k�⦻���l�vG�VF��0ț��gu1�^��0%BR��W<ؿ6�ݢ!��OM��L���J�)΀�.V���������A�'�� 9� ʇu��!��\Z�Z�'N�.�$p�遧��Mmq��}��U��"��i�֜_2�6�ܓ�x�,���C��?���U���������V��Y�2�K<��NM ?���.\g���7��R�Q��v��h��呭���Z$ֿ����un��[W���@��T�q�|���-��=k)�C*�|���")�G��Y���9�3n��z�$x���D�o�\�]e��fQ\L�g.�}���(�������k6A��R�ǝ� ��ϭ�$���hVu�&��V�#�	��A=yh��`�C�/а�����o&��-�!��b2�Ȱd�x�.!hJ���o�ı~���nL�hg����sQ���O�k)�j���>\�b�lki
+K�٫~L/��2T���=��Ǘ2����ug�Х��6-q�� go^��A��@/����q�9�2_���f�Ӳ�� �ji��u��v3�=���J���Np�����-c6�K3�_t����R��-�c�����7FU���Eh��K:��G4זS,F����DE:�a�3a�#74��}�b&qR�N82�š ����?D�wR�&g��-;;C���p�e�h�2vgg�V�"l�>Ss���s�S�r�y�K� ��:B�����R�ps�Z������!��_ݽQmQ*����u�����Qoc�J�e"�(k�d%���r�����Z[[3x�������r4쮞��D��S���I<[�e�d�1���������SD1l�LΌ}�
�|c�d��˗��Zz����	?�r�<׸�/o^��c�r�F���f@`�Bg�$*�[>#e{�,��"��U��Q�#�5��"�5Z@˓ �`�k㘽%�NБą�cS��N��[��4��|����>X\{7�D;%��8W4?������/���B@�psC�A}��7�������"�N����_I"x�yP�>��!1�������ڻ}JN�؟�ڐo:S#�u<�ӈ�h�ϵvv;�L}�Bծ�66B���k�4P$~�E+zM����9�2�f���pX�CW���V���q�����gX�����NEnw����90^��1�2P-�x����Q�8H��ژ):������bǉ��;sw�^"a��ʨ�Xm���-ʳ~� �GB���.���d/�)|��I��w�}h�gr�g�KF��;��=��t�v��ţ4�W����DI�B��,jN��B��Y��Lmv���kd�=�W��T<C"���/���@�# -�y8���1su���t7R�8�+�����{W������,�,��H'�:ﷻ��w.\��m%�a�T����g��n��1{�f�{I��v�7�^���}^�z|*& �t$����hko�;����bἎ�����Z^�c�,������f�'��� �*�7,�d��)�!��$�@b�j�hp��L{�#Xkldw3���$�..^W�C��L��e�S4�h���	�����{�>4�gS|�SN�M�{W�ۯ�[z,�[��8M�a���>���2�si��F��.v���T�5����$V�k��a�G�=[���͍��B���V����V!G�W�؛��e�a|�!�X6!l�����}�"���!�hgWU�M��L�-:��F���>�0���t�2��~ReEA��|��C�w������:��!+�qރ]6Q���Jn-:�2:�1��xa����5xm�R�R���_�/ϕ����St��W.��G���֭r�_�quD��u���`)/�A�����ۘa)�I���������i<��q���
��e>i��rvs]�P񥺷L���(�:����3��B.�������T��ܒ�	������0�����`�~�˼�S4dG�5�!��f�b�{��ƈi�r�?B�ܳ��6_����4�{r��;,.r�sw�I�K=OѦCb��E$(�&�GT�Æ+n!�dF%'�ߋ6�L�<���gӬ�ޟPUR����򰯷^�G��I��1�<���a�X��>$g����rww�o'����SV��½nlM�~I��_�5*&��9m'�{��C��|~#I4V�'P|�J�G�'Bū*�&'��͞�ݱ�,����%��G--�Uv��PL�~B���a%�&�� �,A �h�EԷ���h_g�MKT�ط�:������`)����Q��l�b�k��HdT�+1@|��~��"��c�}(�S5�����ڷ��>�n�\�7�� �HI�G��{���ú�SJ�'u���gJ�.а�����VZs�Ke�)�/�S�x�_�s�ׯ�~��c�pcL�ٺ�\�:���!��%�ʋQ�@ޯ(+�����V�<�����V���f#����귡Ǹ�l�nlX�l��lᴗ�Ƿ��BB�����{"X_��X�T/'����Q��DW) �O@��H�4�^�0`�h 
�^Gou�P�6�߾�@�9f�[ў��(Híp�&���xt2�b�>Nrņ�`�������m�k+"`h:�g��{����)^��w���w:
^B��?�0�M��K��0M���r����z#�)���ڢ
�z����c7@*a(�� ��K�A!Jȴ��x�W��w��M�}�ABѻKP�C�r�������*�{���5Ӂ�J������ی���"V��;?6^^.�$��;vgz��X�/I ƣ� ����Ԑ�f��q7|�|jRy.P��}[�{/r���(�p�];�ܓ6$�	q"gK3,<T�0����7�;0m�u��_�
�ȇ/",����N�l0�0:k����;q\Ee;��1cotɩ�L'���[��.I�8o��j�݀���#��� �h��i��@-���y�>K�}g�D}��Yʟ>\LZ��"��/�;T��ϊ.ERC��&r�M�-Z����O\���uAc�c��:�U�fNО �jɔ�W�P�~7��������++� {��gS�ѥ��s'S�hX7q�s�ѷc6D߲��(�뭇��A�Q`*�Ok^����.�����!O��2b����<�)��U��X��#����|��|��e�@k�C���ڏW�C��X�/���ΎM����`f'BB{{�Gg��]at��qk�.؉}��~pX��q�s��B�] M&��Zo��;B�[0�Z�\;�nDo�#���E4��T�Z!� zS5� (W����ݽ1�{s�
p������_���yQ���;�1Ҫ�fqM��3|��+y��c�fs������NMc&;On��_	B>��sc7�T�VJ/�5����zD��f[yw/I�����9dd}S]/1^�t��8������g��6?�1���8�b�?�2�Fp�l�V�$*JI?��SW>�@ݶ1^��~O���q~c�Px ��ʲR&HT�GN����vbS�8~�^��qBH�qr3Il�B(��"���޲��u�w#���mO�E�P��� �å)P ����׃�?VgR/�j����d��`�/����Fr.cC�3�d�V��~��}���/�8��=P��g�qQ��k`f���<�Fw�1@.������m���  �<��'y;#��k��.�L�����U̵�UضC�t�v�_/�j�XTG+�c���^4���ͮ8-��o�� ��ST�y7(i��̇r!�R ;A@�E$���w��W[)��^����9�f��Þc�,,~�߬G)�>h�yO����A���-+��D	ģC9�l�9��!���/�V�I�vq⦩��$ߥ_�ŕ�fT�-�R֔iJJ���M-lP�@�AF�M/IU�[/����ҡ����M4x�\U�x:_�&c��6�+	���VX-��<�厅A�����ֳm|&L}4h���0����ȿ�7@����.�~�0z��ɸ�-��}�#��S�k!D���U�A�G�^��$D{_���W���<Xm�=d_����YsYQHdx����v�&�<���1mX3�=r�'ԍ�������@��@�=,O�����`��l��&[��7��\�����+�����M��X��k������W#���ND�{��O��P����7&DO���p9�������M�"���$Cy�o�m�Rubw*�f����O�Rn����z�nY�-���&w9�A�3�r��_�<�gf��Ty�"�=n!�N�Q=��d�:2�����5[��9I���Z�&����h� į6�s�M�:`!v��� ��{Yr|v�#'�pq}�E
7��3�z��tE���^x	�L2�~�,���k��Z3Q�(�����->�,[�0���,��Ib�׭jq��yvb�,��
�rkX�r�x#���z���e�jKɉ��l>)Qd$��~�]�rp�	dd}�s4d#�Oe��`)A�@'��t��B%K��d��������,N���e����%��ϴ�O3(�~��Bm��ײ[������ʏ���5Y�x�J��=�9<��sk�h�9�)Sx5�7{�C�9�]�ő 'NS��O.�g�/Ц~F��i�2��%���Upv^C� ;���a�k�
��6C[����}���od^|=��m)_-G�[���ԍ��Y��� �7~Y�vNտ�mՀ��X���cW����
�L���Y����FR1���b��b�q+C�?k>�$q�������4��si�E'��g�t�q�:*��8/��vYEMU_ki]a19��6�JW�b0:���b��w�S����;�!٪�9�ا�$C��Y��1P��L
�� �fd�VI��7^!�t`pc���!�jf*������WjOS�7��|7���ķu��2�� }����qMg% 9���4BZ�
������+~SD������k51D�4��W���&Uo�Z�K�;U��4�^_�C��=%I�]���9��5�OO �N�X�A����y�y�[�=�B��E�'�|5���J����O�u
uN��l]\��Y�p�܆�~)�W���C����;g�?�d����Ӥ��o�1�����qۏM��ͣ!�mϵ?ݢ�c�e���յ
HT"��*�B���Q���FJ-�ӵ1�N��#��� fc�?�(�9��ΐ��2Z� �,αςxˍ���2̽E�|�0 ��D��`�1j�Z�y���Į���=O`�seU��ҫ�:`�O�^SZP� ��Ce~�W쵹��`���M�����M���\o	^�'u��#M��p��ó�%�?��W���3^�SL��~���Ϋza$�d��zv�ʪ�X��^g�*/��$� kv�#s��"{����Jѻ���I�Wº1�3�d����x�U�w��*.|��Bճ�����	��e�7"��G��q��wK��b^�y�g�1^9r3r�?����QϿ7���N���R��Ԕh(2w�\+�Μ�l>�OI��a�wY�?U�;�R4ZΝw����ү�;����^w~��j����ZS!5�;�k���Ǣ���&.�6�P6�+�
|���:ZY�w��&��zج����MT�mrn��Y����?7M����E�M�/��~K"~X��8�"mx������k*g��~�~+�����^*m�#��,�pc3x�抓?��\��(KC:2L�\�"ٗ�&	�x��_��'�5�͈�_�ըB�㊘l�W�wg�BܰI(����Z���t�;��I��~�W.�Jb r`���JQ��H��^#�����A�ǻ����%\�'ܾ�,��b�6U.��uD�ǝ�g,!�G:ӓ�/���.��se/11Zǃ�1Tw�F~uPy:��H��9�;m�{#�����w��cc���(�je9�����Ɋ(�~{bh��1�3,1�(�N��d�JV�#伎;��i��@�
��M��c�`9���8�ٌ�*�.m�}���I��*��P�~��q2gex����l���������C�\�!��x� Xp�� E�Sp����q�����Z9���&�hW�_7�.&.���`揁��&�/%,^|��"���Ûw8��!�Dԭ�Ж��Ϣ �f��:��w��/�Y�
0��>�%���@�F�W��|w0Sto��bd����U�Qb�������N���F{B�����4D�6�"�੶�ٓ�"�W�Z�m���b�޸�v挿��w�����E9@�n��9�͔�A[8
r��&��fdl��I�Z��Z�5�Z��jj��*{�ε��am�^��H<*�Ύ[-NT�F}]U#;���2� C����(�]�z�@�W�[��MPT$�9��1��
s��1�i����?���w�� �J^��Օ��9��۔�:����%�2���C��F�d~=����QF�FE'- ҉�2��&nw3(�����P,Ρ'��Z�v��%���/�F:!3�B���]^���l� -�002H)
�Fs�IՁ7�6���AA��ͥt�M&�z��g�L¶$�����σ��Y�m�I��%?�t�ߕ�זFG���'����Z1s�
Q׈s��Ÿz�n��+"�W�E*�uSN�1���S�>���X���gѬ2���_��=Y��τe"�W�����G�p�Y��]�����I)Nr�:S�(g'�7����I��v����)���y��E����nN�pZ��?�D)���kخ��p4:���TZ�'!�3)^s
���z�(��H�$;������4ڊ;mȁaͥDR3��a�\����yU�=4�	�_�;��I���EUb�����ԏ������#��p3�0ȹ��0��������O#-֠��`	V_Ԅ@Ehv =6�:�f��p�9W�ܑә���o�s���G"��ɨ[�_V�^�3���q�^ܜ���ZZ�RWzzB:o=���o��3��=��s�6r&[��	_J���vu%�_�!���x)3��,����Ah��J܊�L�)-��+�p���'�}i�:� ~��0Qd0u��<SK�_�Z��SA�[.������[�"y/K�����̷ii#�vӐ�e"V��U�!j�b�)���2]��~��=K�tE�����U_Nܗ����o ��_L"�jUkV�)����P�D1����=�_�	��$��Rm���<X[[���ʔ��9��'\�z���S����z|+CU�S�o~iS3��ia�O�p��V^��B��x]�(����)��ʏP���z�q��[���+�}D5#�v������Y�T;�K0��-'�2�l+��̻!P%)�oDP�{B��҂i���ɗ�"?Z*I����ň�u����E��:�-�@��C	�H�:�,���D�1��s%�y�l0�|��o��<�%����9w�y�B��I{z����J�o�[�<hg���"|Cq��Zr�f��~ZQ��� $�nĮ�� �m�������[$�MEQ�^��6?�}�o�I�aW�۰<T�`Q�ݭ����M�L��p�2����ͬ�	-ނ[7UQ�v�-��\nߔ;�5�W��a��`a�8�PL0���y���ֳb�5"3���(=崋uc��`qL�*�	Οͺl�p�Q�6*�́�lqq9)��JE�y���ZX�0
 =�xB�:$�ĝ�xyy8㰙/..�/&D��Ue��nS�{��O�Ue�/m
ѾW��ͳv0\�\d��?�4A&�^�k�9l���g��I�y�3φ�����CT,,,%�U�ԕ�n�>JV0�ݳ�n���e:�Eʽ�=���0X�_�f}��g�yߖ{9ݎ<v�]<�����Ł6�0ʌ��7v�W��Ύ
�㙆�+���F�@ddwǦ������tj����%�!ؗ����e�,�ɓ�W+�{��lx���ht/��J��~8�	�_�ۜ��60���{�2?n>q�7�w�wR>��D���?}�|D`�?o:�=����{A���9�t�յ�h����"�;9�%D4ז����Yu�?S|\2Y�Ũ]��y�ͻ�*1ۂ&)9������[��h��]��|9hf߱v�Mf�8�[����l�Լ2G��S�P���NEe�j���׀KVl�x�`i�#O�@ET�;-���L�f��֛2���3����l�B���v�m�_�	����y�'��o��}��P���&�Awy����qj~���M��������m�{�����׳G|{.|+Z��j�4��ןx��>\�Fx��A,:�#���>e��v"��n�FvW�ju)*��K��& ���`��S�k���zy���$Ņ��ԕ���ӱ��k��=!�h--~2x2�Z5'h����V�kgGO�|�M �t���X�d�,��Tu�����9+N�����c���,�����h��g�2�i�`	sc-�N}���\��=xk-bo��BY����*�M۵�j�uN �]y���o�В��L�����-�i�]U�/�`.�}K��gR�\�Yk���7_�����k�Zy2�X���04��.`o1��ϭ��.�.V�t㵌W�hQ���8\S,QA�*n�3�.�)���b�+`��Y`��A���~�ҫ�G���Q��ˋH�ڧ��Nf��\pw�v�őd]Մ&Z�Uqd�^'����t�^7��¼mg�q�������������ü�l���-<�F�/n��&�{�B�Ы����Ij[�����~F�7u�T���a�d��B����`N��4��6���'�oϴ>������A冐�~�<p���w �ͼ���,��zaŹ!#u� Pc��	:��n`�?�,��6]Q��F����^x�Z,׺Y�+�E��/��N+�;4��T��B�X�T �*���􌚨G��UDp�5f�7�|Q;s�<���a������W�$F�q��7�4�@7��" �h���*:�<wa�G���۶�k���=,؂Q�}�WL�hp������a0"���y�߭�r���7A���e:�5��$�~�����*��Z���=�K����(�g^����l����wD>�x�Y��l�6�k]��B�:��α��u�7�<�VF*63Mb���n��B�m�%i��f�BEz��	���� �ls>#X� �.q�Ր�)�ul�kʴH�s���Q�A�&H0��;���=:��m�pQ:�����^?t���޷�N<V�l^�k����EXٺ��;.�o��zYwƝ�0Ư���DK&
.{R�V0������b�ܳ�N�׻�{���b��v�G�Y�B7k����9���/���^�	��ԉ���os�����0����%��Q)�vF�/��wY�&��WlXu3�}8%a����ž,�?��uŹj�*�'lN�.�U�,zKֺ}y�ݵ�?��<(v[IjRc��a�+dY���	h]m f���m�g�^��?���-�Q�uL�yBb��޹���O/�����&#|�V��=�hb�ǡaK�g�ӎ�Cay�p�O��Mg�Zb2�n���}o��69h�����P�S�lFlk�򿾕�8ϯ�8�5W��d��-�<�U�����]t����"���yȨ�^�txx|�?�c��p���Fق���ך�Sކ`�E��:0O�����j<M�u%1)�"S_<P{7�O�\������q%�aI+��<A@�0q�ҧ��W��a1|}���C^z����uB9N2����Y�əq4Y�((�54�>�B��l��l�se8���L�x��+'RZ{�		�Fp-��|��/��?\*y|�A+̅��GQ{����"���'r{%�zX�6��#x�E�c��J.���@�[���
���}0��-7��T�Yj}-A�CNg�NX��샩�%U��X���ȣ���]�[;���x$/F�BP�?-��4������v�����5�y�C�nw�kg7�0� 8\%���	�+Q�W-B*������͙�a��G��ԛ��!���=_M�h|h���lĐ�=T��Z�ج~t��sJ��D.���S�_��:<��E��wO�����uU��0b/3���+�FN*��M@�_��|4��o�����l���2ȱ��\�}�kE��	Z_�k�{;��3ӿ2F���%���Q�C�n�/ևH�!�26�{������Sù�	a��j�w�T����Pi[q����45����i���Ј𝋑Y��2;v��moo/���s	ƖT�E*��r@\^�a��kF���b�K&������{	�o��}��ct��&�g�-��1=f����וUj����y��� ��u�	y�wp �(�/9�\R�������l��ԅ��X��B��k�Z'r�8��Ki)1��e�7��+���ѯ�>vh�����Ha��ϋ���$ߧ�ׁ�K�V���r��Uч���/(~ⴇw��Ŭ�����@0z������w��k_o;�&�<8�i�����?6H.�L�_���򪱴��e���M��?�Wr�S_f��� !K�	���㙁۲�,��,���ѢơL�'����e��Z��0��|�	�(���5�F����-��j
Paܵ����r�^�x��������=�U_�������y���M���ECx_��к�]鉼ԃD�e����o��W ���[�0��Z�I4X�b�WJ���t岱��}�%m5E	/�
��m,�� ��jֺM#tG��������&J�K����� �����ɵ!/uQU+�J�Û��l���S��O�<�I>Y�O��{�छ�<��O����=X�g�7;Sl$s��Zd)z� Ia��ݢ���=ڸreE�~x�Ǝ,��$Ҡ?R��q�}���1��=?�x��6,?
0#�h�lԸ��y��
��R=���8'i�Ǔ	�W�]��7Ҧ�Lr�t�\�|���;3.���1ki�E�F���-��O��J�*O)ahe�G�\-�,�6��51��S�Ŝ���f����9�b��D����ﲔ�~j�=���^��9i��f�~���}�a��K	`���	5!�����-�{��vU�R�*H��M#w��C�i��P�)i��ςDRqh��dm�R�7��'��rOk�����o��,��o�&���3���v�Z6�B"ǔ�F��I�/>S'�����n�a��Z�q�����|��x墅�ؙqx�叠�Rh*�NQm-&���eF���6��z0*�QO��;��[�f�����o�מ
zi|�|����1lƳ���|���[Oi<�4���v�GYd��'��'�:�xc�H���݅��*�^�iS���
��:�h���9$����wdN�Jg���Z�����Bx݃��Lm8�~c��v/<���X��O ��7nUī��\��$��*���ϲL�M���b+�Du������m6�Ҋ\v�^��s#��)�45&,��8�*T0���*N6Q�k�YM4����{T�����h
��\n��pJW=5���4��C����Q�����Pi��$Gǐ�n��nD:��F7��g|�����{;�9��9�:�h<��� ��z2ֽ�����������/��z4�� �&�۲�@�$���D���]4')�0����x�Ym7=�E�
p �.����/��^������8��WSߐQB�,ꛖF�D ������zM��b��/K���;>(W���N��-��������d>1s�R���lIŐ��.9�Zo�	)AHh���h��<�	�c4�TΤ�7�7z�����)>��z���[,�npN��O"�Q���T;l4�<�c���k|���|��Q�[)��QpDI��Gţ��%b�3�y��e@/��������;;g9:�k9�D5XƝ;D��@��5oi���
���^����:�6�r�QZ�܊����L��7 ���V�V�.�&]�{J�s�2$��ʊQ�n��8Q����ߗ��=���F���/%���Zjyw(h�p�PV� tƙ:�p-V��o�� �"t{�k՜��ly���T�n��y '�R���u��!�I��.��d@��hY;������ew��T��ڏ��
��Ga���������{4�I��׊Ȧ�}�(

hi�%�o��N�6q��ݻd��G����2��/�'�^K~�"E��LU�� _j|�X����$�<��K��߻S���6cUa;2�4�#��{~�$�Y�?B6��v�G˅���^h���!����7�&D���"�_qYK�}B�ҟ8Ű��I$Y�z3�W���~�1��4��	�$�M%���e>���8����{Kfw�LR��������ߝ_;��Sk�����'��ӳk'�1WlLQ��l��`"�O��m���RHY\Γ���ۼDZZ�9U�[�Tz��p:WO��ܸ]�<��7]N;?�����GA����x���(������H�y��Sx��nw�S�Ŏۈ�p!�C4I�(��q���Ɵ�	P��.� d�$1����B�����^j3�	��9K	Q��<�=:X��ځ����������.���֪]V�cum�ϋjG����Z-ٮ����Ӷ;�P�PiP�<S6"ȣ��(0J1Sˋ�=.Dpn�譡l�>ja���3��m2�dJnL�[h��G�yӯ0u����x�,H_�ҭ��;����x�);W^
�T:�H��~��%�~�U��.�h��Y���ɍ8�|���%_h�P0��a�Ƹ3��!�Ci��b��ۜ��.1��@�����4�]R*�o��$�H�T����p��*o�x�)��}`7�������㾵��6u����@���j\����d׏C��QZ�n�/VO�ev�t�h�b� �w�I�9����+����:�j�*�Ep@��4��N�	�7RL[�z��x���)��FQ�č�8�|�P��S,D��m��m���q��ɥ���䢞�X[���� @�mB:}��[���y���N.�/���P�����3���'v�qye�����щ%h��V00�Zu���g���_kC�̱���
��{ ��������n�����'��g]�M\[����O7J�CI�nF1;�rQ�U?��9�S�������4q�����^��B��dyy?S���G�t2�:(�	�+�[꘣�+7�FtfgHri��j��]m�[ I)��9>���aJ8�����B�b��@�
$�G*r��L�ˌJ��S����}?�0����sc퀧�ߣt� ["�L8Ե�`c� v�.�H��@6�5��m��v�}�����y&�8�d�}*S�=�7�1+7�2�p��?u�=��V������1����\���P7�RHvo�+I)��~%�|؅�M�%;M�Oqnɬ�}36g��׳�����a��+�ԫQal��a���$b �9ݻ���6�
�3bn��\��:�G}�m,�u��܏)L��bQph9����y��4�
����AR��yR�b�O�\���,���6�իv\�r�=�=y�/N��f$�z�]D۝U����D_�����sZ��E�M����0ϡFg�N�#�����ԏ�[��$��,���1���?*��U%��>���e2��7�����S>�6\n''|�c�l�A��z���w>�x�{6�s�dax#��V	� �����M?��FyQC*1 tb�Պl���h�<6Jz�im�񑟷y��%
��؍q��H֌�����Oٛ�vE)�6��"�\5 G����y�T�1�/9���J�2�!7�}���2��Ä&�qU�΀,��&IdT`�����Q9~�xXZ^'���ީJ��R�25MX,͎��1�:�c��~%�995��°���Li.�F���{���Tp|ݪXc�7�,8b�b�Ѕ�UȤ.�s5�!b0S�� Y�w�<2af���)�HPET9sP�5�7m~(o6�K�@�m�#Bû|*�RIQt�<)�|�Q�:P[�A�3C0�&~й��?�>��͵����U�%��w�f�i����-Q���<�=Be�{�_����:Z�m�*N�{F�����V�&*�/{Ѯp��)��M������ٺ~-g�����[�V�ǿ�� ��ڟ:��w���DU�ǻ�ǗY~b�.vr� ��	915[P��Ɨ۽R�Ao�I_�-�t�sQ��O�*o��������D��16ܶovVôԤ��Qy�%bN�8���y!غ[���ѽ��I�+���.9�_������qE�rA����?3�j<~�3DAe^zڳ��-|�W@�(YR��xu$Ő�"���.�z��[0!/t#lc_��F6
�2���r�~}��t��P_�ZB�r���s>��j?��c��WtD�
 �G��Y��peN��ii)�PA ��&�[�p���T�M�
�Q��^s��}`��H%�d���f|��F�:�ܩO�T�e��ٶm�N�h�.�F���v<��ll�V�k'ӭhDf�Z1P�aZtX�	���ǝX�'Ϣ�KQ�f����0Ƨ�ُX��ߩ��}�w���ƺ��!:�t	"��2�Zw�G�=~X�ܜ��j-��{wQ��Ȇ�"��תj�ܞ��|cm�9�Zz4���!��i����[AIH�Ц&2� dD�n�U�_̪�Irg&�3�H�Q�)f�=��?�L�̟��6��
���ȤDϞ �����8����Pp�N��T�椧w��d,�;B[g�s��#�5���V^�� �K]G����r������#�o�Qj�.y3�N���w�鐹z��S�� aV�R�_���b>�eG��������Ʀ�Zo��D���Z_�Hmb�k�39�[��Uv[�����

�K�&$��?ݭj�K��3z�����4sXUh��a�����-�k!J-��zQg��k1�p��`Y�ͰM|$at����XH� {g��%r�h{��FX�C����}����h�`�L���IJ���WJ�
M)��7s��̿[Z,���}�-1yg���S}��g�0 /�H�*�R�RȍH��'�ZU�9# ����X��'�b�ym�NA+�P�)���`��?�zh?���{��8�����Lwq��6�O��$n~X���|\[Ӕkn��=4�?$�\� 8iE�шY��ƄtcB��}6����%�����Xi�L�D�0�3�M�D/ϼ�F�-��f����b��.�7�\�

�N���3��&�D� �D����HBq�B/��S����3W�����+�s�}�]L����*B���Y�o���w���:E���Rk����l-B��O8H��H��Jpv�y=�&��S!��"*)��':��2����kW��	2p������c�[��m�yS��r��Iu�GO2�VC�h{K��Pip�p�t�J]ڱ����vr߼
�1{s�@�X�ԡ�����#��)�3d~s�B[9ݎb..�L&�<j�|؉0O�۫:#��Ol;Hx���(���j�_�ڪ�8��U�̃K:N����h�B�~uy0���w�nG��E�U���_����l'��(�X" �ұ ��k{�q���}�U�ᩛ��SSS��<����@i�:���μA��G��<E�ؘ/�sM"�����Tr-�i'L��?�'4��R�3�y�.���a�_y���6���&��JR�h��� gb�\����-:-���V��������r��eZ�#���0oT9��#�����ѵ[X �o�_|F9!a���|����<{��xĖ��䊹�����;@�@�LJ*��.�6Ń�)5b.o�-_�=���W�״�i�x:713e��Sѥ�X�5�s��1~�\R����5���n��E)4^o���;�c�:ZL.���r�ςikk�Ꭹ��i���V�c����trt�ˡ#����lua=�����%�"r�x��\Ѭ����u1����e-9��Cm��(侲e9�ޚ��O���4��<܎��@_�����k�#!;#ؘ�o%�^@�*��]&��KO<��8qi"'UY�zS>�d�u�la�_�����<8���׶v�x
	tM3�+(I�;sѶ�)Ô���P�@���{�]�(gYk����h�	dſ|�O�|g|I��s�����:06_'�_5Dqs�d<G������ʗtB��ۯ�Bt�̄s����.���,��͆'=$��Cj븗��b?�Ln�u�{�|�2��b�m���$���;85ϩ��'���PM��L5��I��?Ύv_K�w�m�]�7������#n}=e��p������6�"�F\���B#�"C���^��!K�SK��Pf�"�%7A��Mt��
�n���1���ƶv�=!Ƹ
��c7�W�X�yq.��M����Ìٯ}��3����i���Ѣ�z�XBؽ��|�?�������lA)��(I����vS(H�e�J�rL�y}>q7�VJ�-��1^�
G�-���V:,����
�iqs���|ԑ5��da9g)_��.#b{��4=��������{�	��6�ȅ�����D���(�3�"������223&�4�@HS�2�����Bv�M]Cչ	��Djs2�Z�s�]�Q9�j�9vFT	�<X�Ŷ�����0���c,S�A��T���72U�Oa^p'Ml:��������*�����Dp��pI�"i6�)e���@��˯���&��8�p4�^]5���xo�F���tp���\?|r���D���V�s}K����z�GP����~Ҝ�(��=��5���Z����<��/��g ���I6��h�s���כ�6ܲ�o�ݯ����qT>���C+�u%Y9���)�Q˛��=5u���E"���[P�_҄;52��F��>�:��!c <��*����hLK�>QE������;��y��W+~�
��O.<c�ݏ�wj�n-��{(����^ݷf��'c�ZBQ�T@���r{%m撥�MՓ��ذ�ھ�#��y.j�C��5�vA�b$���m~$�4K�T�>X@U��N��d��w�}n)��{��/�>���.��*%/$7y�)�{֛��#�D�r|�K���I����5݋�9�.qp� �է@�KzO�>-I�ܠ&�H����S�y�ܰ��!"@7_/�MMO���oPe-�]!0mZ��ir�6"3��X4�#/�AU�v��l�&PF�=}�9�=b��~�ϙ���LM.��ۣG��##�5�Տ�,T�� rh�)X���p�����5s���\�÷F�
;:���Q��2ܬ�열��~,� �v:g����\�>�ᠷ:��V/�O�p��"�yil�X�Y��Di�~�\�j6���&�R�Oyi������m!v�]�*;���0�Kq� P���[n��EV�Sc��b�ge��V�`1�r�	љ^V$K���#��f?�7`p�cI}��[:S(�%���1G!�D��%����j�����綧��Oq�H���1��m��~����Rh��d���p�{��Q�7��7��n�c�o�wdJ��Rmh�w3^�:�:���jF����)����P޶-7��P٣0��#踀���z�$���P��-f����\O�G0�#��JYA����]h���f�S7�Hi|���Y�>\�p�-N�����b�ddأ�d����2�A��:��/��vM^	>�Rj�b��Ge�e��u;m_���;�`�*�@�[<��3%�]Y)4N.����uz�#����ww=�XRKl~��6�q};��k���.��y�[���ΑG�=�7z}�=	�E��;w�CXd�r ]$����W�T���E˺3��}}�Ȇ$��n��Zͫ5Z����t��,�=#��sMaX�>drZ��~E��jp*j��
�Зu~6h�߷�[;�%&!y���QB�-�ɫ'8P����M�ҝe&U��MR[:���
�b�5����*QbO.`I~{�t�bY:�na�ǘ{�]}���J�U{��M�- 1R2����G��_�jA?���X��U��t`Wbh�v�S@��҃է�����nՒ'oH���nv�}w� &���g'r`��x��z�eN��}~�^�\?<Oq� �#���bgM�AAv��6s���I���]�'x�������R��!�(�W�*�"]�	S��8�~K�%��5y�GAMT��s�(f���͎�ܦ):���9�{���~�׮���[�G0s��G[%G[%�����់l��,�iYqW�+�p�#�g�1%��y�`�P$P�d�s�ģ�Wn��4-$��^�	4bE�>\b>�U��/�Mhhg[A:�o��0���hWz[�����*��9w�]���]������VÆ�Rj;Se���(�Lz��?���҉d�/8��(�&�j`�~`΋+����rnG�u���}���~衃i�>`X`��m6<��;���N��h�MmZ~�����Υ�h()O�]y3�rVo�p�C�	b�>I�z.f@=���ԩ���t2ep�*̐7ò�K��h�R+�\��[�ݝ���%��b�Ä�y������=����~�ط�����.!�C|���r\�x���zp�72`6���/~I6rJ�������&�i}����)��:�C�Qs�W��[I+�7�`�_1��A�?رJrn��.�{Zr���<����Hc�D���׻7�cUĝ	ɳ��͍�*0����w�U����rm=o�8���?���~s��,����}�;�W�6�s-�'�.A��!l��m�s�y�ؗ�L�7�l�\I�ѝ,w�kF�`o��mh��Ѷ5,R�x�D�wi���m�Z�=b�#6�v��j ����{k���$e���k��kV������B��ŁNL<��+$���D����1qWK3�V�,�L8�߅(��m�(�/`�IZ�P�ƙ����̒��I����8��v}Ӂ-�*��
8�9�٪�{"����nU�w�2ЍC<4GD�(���J�i��j��<J��o��ٙ5�@��.c4�_���v,x�~�����ۙ��R�����鹺�	�����	�tAH�P<I�u c!Z���D"�LYQhH����I��@+RZ2V��z���J�����蝚�ob�-w�T��8O�y���|��=a���͹��?��d?� �М�<({��F�_`��u���#��(�V��g-%�z������j�y�-�;
2Z�p�M������a^Ͼ���T:�3�����r;_���':�U��"iW�+N�ΉA��lƚƨ	�z� @M��Q����81h���_�ܣ
��y�Ϋ��1�`�>�� %q�Ƙ�����p���d�a˭�K��Ki�7ۣ�&=�5�jƒ�d	��wzS�����	�?Yv����z�E�f���0G�[x�H3���}���q�+��Zq�	U�*C���f<�{S�3�au�&�l&�⇒`/'�@�:���q�A���|�K	�H�D=4J���^PT�Y`��D�O���{}���of�Aj��*ڇb�ڹ<��������Gҝ��U�:��@�>������FLە���V�d����8��GKf6�5���<F5� eBN��;{rW s���4x&~/F�)b*N|���M���p� ?g�o�F���糮�J1ny��ȕ
�K�h4J��n}Hm��:��2���S^ac�!�{q�B��#��,;so�'Q� ���5B����`��/���������6��|#���2�՜
�;o
���|�[��xF���К��A:?�EI�������)�q��ũ���$W�~Ŭ���̐R.�$�:~�p~�\שa-N�[�7���;
�U���w�pU�O�7�H*`��9��Z�a#�v��D�6,u�v�i�f��y����y�[U�yUr����y�_��?�VɆ�Θw�]l4�0#�12|ii���k�l�p�!h�)a�m�^
tB#�Z搪�1��X'M���;ݘ���0����˞P�<X�Q;4G9������ N5�h̽�q�R�;Wr��~wT²����̅��q.�f5����b7��-O�)�x_�iMn�zA}��@�Hr����r�*c�3����f��sH��`�2(w��9�������;��ђa�f��u���F��<y��O�K���)�۴JW;�D�|}c.7�M�rn{�b8��,��x����;qI�?;U�&����l�H��MUu�<�E��Z�X�'<����	��I��Z�Y'�r��KmGA��f��8�|^�N��I�0a�Vޤ������u��3�7�P�'����yX}l?���g��[��X��}�t��b�����V�~"�P�AD�V�^N/�Y�(��;�ABۀ�'N�'*�oP�N:pT�W+	���sK�q*���D���Ò��1	��Z��@����ӡ4>ʔz��/
�^���k����|C��nM��8�7����N��?sZ�5����S77�:)#uw"�*�`wڼ�gb�tF}�b৤�Ů)W�Hf�f������.oy����sH�ٕ���*��DI�bRk�@(i\��^DZ�D#r���(_s�f�8Y�:WY�y���qi��A���/��'�6�s�QM!�3�A�vP�W}�AUN��MF���ت_�pQ%�+����|M��M�7��XVU��[)<"����BK�f�G���Ό�Y��w7��y=�5�=˨�p�P��P�|OuyЁ�m������-EW����&���z��9����9HpAV����a�aDޕG��:.s����TJ�ރ��c���Ԙ����� փG����h ���xKZ�.���s�qO�Ϲ�fN]7�#��R��@�J)�s�����:�qh
��:�������\��\�O5E��S2e9:cZ�������	U#h���3Q���T��A����A]�|������#��ű�bf�n������bI _��41���}V�� �_��>v}�K}�6��;kO8{|gDnp�q���Z!E\U͞3�uU��ϙh��)��@i��% A	q/���t��U]7"�#d.%�6Sn��VL1���0D9(m�$CR��s���?��l�u,N��m�=뺈�I���E����/���W�?��|$~�\f�k~va��Q��E
��(�JT����]�&�n�3�9��(#$1��
i�eH��Ǔ�n�v�9�5l���&W��|]0)���n�N>Zo���[lzZ%�./',>$�.F�׬������ߔ�&����s]��ư��tƀ\5�9�P�DK��i�V���R��\.筎M�kX�EV���&$��~3�B~,N�I�~©/�:c�1�6�h"�I�'vU����g��o����x@��tD�*�1I�a��w��R���UE�W*�I�X>Xn��M��PW�N�i�5�<BH�����ߋ�5�6�Ct�U�b'+	e=��d��eB5�,Ӭ�BڈUR��9�}gˇ��
^��`�d��l?��}�\�1�#���Al�q`�/�N�3���Ģ��6�8y@%�@����m#g��Cc��%�����˷������`Y/JI(�Q�f>6��	��͸Uc�\B�\�~p���|x�+���������D�S�(����k
�E�s~�������ZBCS9�@�K;�`���!�Q�_ID&���$n�4�
ۑ�`Ẃ׉��+6�d�͵%��7M���S���� o$?�EC�<�u���N�v�j<o
�V!�t��O�𑆰���Q�>�y.&71)Ϥ�BU!���=.u-�D��Jo������]� ���ݫe�M�;YI����h�܀�>�lZ�;���X�6c̈���f����yxr��aD$P�z�ʊ��&n���� ��*��Kf������/kA��~��j\�D��^���{���ԌwX�I�\��rF ,�:|��!�1Rٙ����~��Ap���o#�tڲ������߰U?��'����Y^�qI�P���'�2�	`���Ғ>�J*�F��-9�2j�dU��f3=�@t֍9�Ŵ�<�y$�p��jӖ�ܵ\��^g3Y|7B���i_���xJ��h�6����^P���iw�1@�Zs�d���P�͹�G�w��{H�9ʶ����%�M1���_���?�*n�o|� ��,/v�˯��r��\�qU3i5+�5ńo�[*��V�����������-	��)N���#��Ž�n�D��.f��z�<������ϔdIm�a�܄޴O��쫤����o�4qG�Q�J�P&erV��	ei`�&z���M֟9��I��(���f��Hdu�}[�0ź���>4Z%z�l�$bg��gjs@��Y-��ר�g�B	�^o���7.pO�4����@!ta�3�MSj��1�5��j�]�V<2k��:Ǥ��j�?ЌݐK�d.#%���m̃L#:ڕ������[�Iob��{��uP"�[;:~ �%lR��mtq4v^qл�-.a�Tn���d�5e{u�6v��
���|�g�z���\�i����S������ʣ�p���vr�$+wzr��p������r��WM�Y��]~M�-!ǐl���%�?(n�}&#l&���`!D��$�W��S��L��ލ���z���#�,�
<�M{���1�*�p�׏��s���i2<�M�j.�Պ��d�.<����K�̉�nY�Y@�4�BrTת�j�y�1�`ǣ�>�s�D,ICȶ�ф�
���|؆��߈���=Oڏ�]��ZE�K��j%��(~UA:H?94��p��0�We�&�8^�q�֮��� �Q`���%�T�U�$��rt\� ��������ee��]�c��*?˷��*ꎪ�H|
5ܭ�� �oѧ�'u��-�[��N��?p��?6��/��o�~���oG
���6������>׿9�#Pߐ� �Z3��ꥮ-
�Yݟp�@��6��-�/���y���zˏB����%I¹S�Qk��9R1Pp�x('���d{p��N ���=|�[p��l)/ے��K�r�I�{�X�m�H��[��ɼ=�P�M�<�����h����4RQ�\����SE��-'����7�tl �:VCx���s�0�o4���~Q�+.�(�u�h���+��2/����eP�7zʤ���:�y�C�x�ɾ��al�[�^q$>�+�$��ƳԎb�}Wo��^�&�#,yL7�|Q��1��>'�R���&��/d-��e��ݞS���;��ށ��Լ?�K�^p��Up��ņ���AՉFآ�L��7ZU�,�������=WU�&p)ɜ�p�	�V���cH>P2m�>�^{�P��.�}�{%�M��{ji?������tUx�]� ���	��:7��!��jIT=��0,[}��>�W|:L����1�)�˽%� Jx('ח@GI½������Z$���͛ܜJ��<JY�Π/º����@��ӑ� %�����Q�G]a�B��R�C���&��"�咑F�����딮kT_���D(��=��H~FE��� �5�5�lt&K�M��j��]=��M4��$�N<v��^�)����LG4�	��]5K���m��d�~��:�;D���u�W�Qȍ� 1=��xL\'��e�j>F3��|�&�Ξ����xm���(����H�'����*��v[N�X,���7����C��T{������T2ސ���D_D�ꃁ܏��}?|�6�M±��~�X��i�Y]يԂ�=��FN�]���s��R��R}B3��^�'�eJ=��n�����2��_Q[���S8�֓�%_H�{M��o%�2tAa�F�^�rP6c��h��> ��������7f��p�-�Hxc|�/Sb̢f>�|r�����:���x�|!��cK�]R��d�_KD�)K��r���/P���zGߓs�؄��ȇ݊l� �҄���@�çU�V��&e~�*Nk�3��ӝl�(�O�A����~��7>���~k�_���&����	��GX��1��-��Ĩ��R�F���O�I7k���)�ږV)'�evt1�{zi�Q<�{!VX�P�ӥ�J��{������iF���O���!�+���V�6tRh���P�!}Jo�8pr)��=�R��Fה����F=���j��5B�t*��|k~�-��-�\=%I�T�"B��'�s��wG�C������۳�.M]�n"���W� �dC�ħ6��͇}��W��\���+�,�lH�����d�v���|"ؒ���Ʃ��n'��*!������Mc�Kzѩ�"eҜ	!Z�KT�{<R|wWf�J�����@��{P��ygCХ�R�>��#���}�lA��l���p"G�;|���W��Ŋ�Q�[W���v��)�ݯ�L)�5��v��gB��d��]y�t���P(4n�\o�8�I��W�|� �9�������p ثӕ�{(87������d�2���.+�0Kq�)�r�|\]r�M}␘vH��q�[��&�"晐�SFq�>�/U)��@W��f?�H�H����(^l���T.{�S+�8K`���b��pr^�dW�lQ;�::<U�?�^ihH�<�@���0�U���R^�bB��M��v�=*^���'���Y�7������� ӭ�6����'G������_$�s��*�v�vs#+�iHm�����a7�X+��2E��-�P�[�����g�����-��e� ����=K����:c�V��r�͔���i���"�A�,۞n�]�f��X����uhd�{�[�#k�2�zD|�4��_�h"��YD˯��9B9]�(�.r�J�{÷6Mg��+�:Yo���3=��z�N��$��2s�0B'O�9[��������%ȁ����*�覦T�̳�?9~�l&�C�0}%Y�C�_��e��<���qgn�δ�O�W�q[oV�$|�1܎��l�H�pa*1^�.}'�&f9�l�eM���
�R^4ԏ�U�.m�3��˫&a�?��Ix�*<��FX�����d�a�.Ȓ;�\�N*�+},0�JGC `{�u�2
gt�[��	��Z��+�T������[����&��@7A;���<P,P�3�ٞ��U=M2� ;V�B�	EK;���n�V��+�C�J;�Y�0� ���$w��"4��g���R����/-Mb�z*������/}Te|ޒr��pVw`"��H��@�%�Z�W����"�Zuז��aOY�:�9u�J��ih(b3��jo���E�ڽm�J
�o���e���b�d�'U�4t���:�U~D�I#�<��MjG��������A�~#-D:(�L�ԾW��ۿn�k�dy��X�j���;EQ�P��/��U�ē�6vŚ��a�^(����)�
�%��A�zm��q�)}�3bF<r��y�9*�����W�6�M��߆$.�*�k_"��"1�MeH8AcOy�BQ�FF�����|�3�bh?`�-[Ce��� ̎T؜˵��Vy��$X��;���3ᇗ�-6�Yw��2�ѓ*�����>�:��)�^	��bs��)4����<uOG8�������/���v�h2�M5��&��7�N��S)l��4�{m���ԣ���]觖3j�� ��s����/���@C�����2�(��n���BC�_[/�M����Z�J��in*% �+�'
��̪'��q{W��,�J~ji:_4zR۟�Jͽ�m�Z��X�QW��JҖ9��d/�u7��u���hj�P�D�l��Iv!$����T����E]̸��/�����2�#�^m2o�?U�q����Zn��=z.���*dODW���;hZ�&�S�H^8?ޔw�-z�$��I�._-/����	<[��'��<�c�e1 ���ͥ0+���<`��0ܖ�U9���б�Ƌ� ���CA�Ï~`��\�f��P �w�'1������ڙ'���w��|�۷���S�A�Φ��|U�e%a2]������hB�w����0����ҹ�^4�*=!��|v�8�k]V$��3��W�$��w9I�x��D�&L�Cl�T갯%e@R�+�����C���y�n�ԌO�h5�s�扶ӳB5�d%3$��8;��M��;�=�x\�+;QR���-�ܜ/˜_�a��\���d�b���%Yo��Qb�q7�Ia䨰Ƅ/N��t6*y���}%8��S�<M][[��&�<�/�Yr.���t4,��uS�>%d�~x����ji��@��������{���՛t�&�C�Ŝ#j��m��h����;�~����'�^\�ݲ&���o��-2C��2�I�Yg�hn����]D��@T�Mp1>��}��#��OĩW%���e*޹���]m�+���T&v@�^0/���]ﲬ��ut�[hN<H㇉��Сd�>�%�՛��i#�_<+ /����Y����B�n�[������}���sz=\�W:ϓy5�$�%��U8���%��Ť������U���k�(��j�ݿ��E���Z���HU�j`�����:|# =5.x��B��.��Sy����l�z��H`�#��b=��x��"DQ��#�Z��s���������8y���[<4>R>��VF0�<Q ws���M�ο��;��k�~���7M�7��T���kΫ���w<����:2�E䧼�h������p����Hź#9��`�vO��P��+�i����p?b��(�`�Em���n(Ky���\�u��ݬ����a� pD�	�՚��'���K��� �}%��r٩:s��e�9��*��9y٣C`<$����*)`n���6i��c��gc�:���_Ȏ��JP%6����[o̗��z����'Z�<(�P���Up��U-�h,�t2�[�~��!�7�Oq��M
���#�@��N�k@}��9�X���
���k�y8�AJ�ʙ՟��óю8���\�}���L]>a{l��^��n����d����Fz`/��ma9��4�?6��A�X�f�B�y�B)��WU,�E����P��6q��|�~_�f�����m�Z��A�Py$�����8˯,*}� :��Yk=J��ҍ��g�����56?׮+�P�����	�~�AȄ��@$]`	���P������-����{"��?�G�i�����Y��ʉ��>JxW[�c�#z�+R�]Ft��\�ͯj��|ZU+ːoO��'*b��}�3������5d�����+���^
�d6cTܪ�8ּ
(,`�		럯� F@Ԫ�,H��hmE���ߺ)#��a+�ǭ�\KZ急�l�����ߏ<��l�M��tՋv��ti�d�(J5��g����t��oy�2��[���^Nh�n��w�>��{�i��+�rDժj��q���j�7t��7�b��-�c�ڧ~
dWV[�_/���sa�����y�ގ� )Q{��*k��q�H�n]s��-R���-��D�x_4�����%��o�t�NS�������`o���;��U �>z,I�J*?�Y�G�W�i�zኺk����Xp�*_C�����b�����	���*��K7"7��f{F��^bI��UI� ��\��S�׍A!�ԉ�!� #GD`�5}�w�L׬ڣ�sy3��� =��o���a���,Io��[� �҉�_A�������T�#�'���z����Aav����SVlM�z��� ^yϿ5��D�V��D�I}?��K����oDu�=ءd����r$�\� 59�(߶T*J��fO��W.�
J��.t҅���У$�1��_����<n��~EC�4��FQ�W=�pzz��j̺>��nK�U!��%��Y�Ω��8�%���˚;l�\�T�>U��H
uÇ���#���É�^?~�y[Ki�WA��Pw�i����f�t C����lF�x�ߞ���h�O�՝���Uo��u�V(Rܡ���C���ŭXq�]�;w�����z��ߝ�g2������k��J�׈r�|{�"��쏞��o��/S�Ѿ�䛊��X���U����A�Po��Y���5H��2%V��3z�B$�l)�����I��;����k��j5�iS�Ǵ�.�ji�j9��▰W�o�:Yk�W:֥n�:X��H;�B�ۈEz���E��&�k5}ҕ"�H<#;��(a�����ޖ�&�D8�6G��9;|_�f�k�_��kS7@$�T k�Hv���t�`�8��w�]�:7쮁a�[����J����\m��r'O�w.�k�Ȩ�P�xՅ�ޫ�����Cwl�~�� m$x�����BHf�e�����:րi��qO����Oz����њq喾�=}���R���5r��#�8�^��e֪��S�Y`�1=��	yeeZZ�9ƹqM�4u��[0�K|�����(��[�<]�(���I�M�G���ѿS�����^�【�g����Ɗ3�Q���]��ߦ7�7��g��l�D-�-��1� t.Z',��2��Պf���/a��ǰ���N9�"4P-��3j�l�v��﷗�j�5�:дE@�Q�?4P_Rx<�>v�����BƸ��L�c�)=x4�$��H�[#����
�g�l���)� �/��{x�Ң;�-Io��q���ז{��v��f�g���1�[��	,�b�@�y����p�E�GR�uV��z|v�ldg�����w�6��P�u��Ϲ�����Zk����ǐ5i��q�=j�^/p��	i>_
���a'�ka��߮aM�?��>�+��d��R��`鮪��6g�;������Xp���|HCwU����c��Lq�ٯ�O�ܛ�6����Չ�T�Ld�YMn��Wޘ�q��r����_��%���<���"hwp��Q�(��BO�_̌}��makh���QTU�c��*T�<������&����LS�KmP<C���=..G���ݮI��L��acC��a�L��f�e�H��XoO[����Ewi����a��~�y �R^��.��b3^��u��@=���_��߆�@��3G�x�)C�d�;<�67�`�����ef[I��6_�X�8��?̖��/���v���.���i�FV�1�0���H�p#D���'xP$�e~s� Yش^���ϻ��_�:����]�1���D�+dx��]����rU3����A%}`��F�u�ju]2P�1�V�ߩX�4�@����������ҝtg�c�,+��N��A�JQ�Z�*�["���u���JUe�;�-#e��-����O����ڭ[H�I81 �,>}nEX#	D�����g��ae���o��Cr*�i�U�~`:���Ӑ1K��hRn�Ms���/�/v�8��,V_t۾"�f���Q�C5Eee�'K�q�h~��7aR�}[�E��#(SUA����5��;����I��UQ�qX1����y�I9�1����[���-~�{�!���7{G�`�1r�^��eD��Ɨf���e�}�J���ʍ�~ͬ�Y�G�o�:-���Ս��6u�lB����3��\1�*sЕ[�-*�����[����_w9��q�{V��^]�xrgC���?p/I�4�Y�����'�,Ci\S�>�%�~���+8q���F���#��#}��so��NH��9O[pD�ƭb㔛��El�(Q�ߜ��f_�)ů-̃3�UȪ916�k�\w@55�/ŪX%�/�L�a�tU.gzx��R7�dɞ',xzl�m_�I��s;���b���U|�[d[�'�6������*8i�:��%�~?�)0l��c�Kog�E5�3i���":�ٴ�d�"�m�ڄ�<ԍc���I�ros��j(6��$���z�����1wl�~��a�j��%l� j�y�m>؏�*2�'�[��~&i��h��y�@��Sӝ~�h���>�W�<�����M[(0�g5�=���6���BX��(ٷ���	�^�o�����I��6I��B϶���T�������vg���,+�,f�����U��y�`Iu��5���c	9�	�nݴ���(��q��M���x�ϙ�u����>`B� ����mUa���_-_xr&��)��eD�S��[&>
����|[��^0Ll�Kh��u�!��k���f玜���(3�q'o!F��Ʒ�'�c��_�t�UK)̙����C����|�»W(�B��u3��V >�	�8d�{	.�U�,Tj���y~��g4�~DJ��'�aȵd�E�N`*v]&ᔙ9�,��U͔g���2'��8�|C�gR׶������ LY2��v��X�N@@Pm9G�y9D�nL�+	S+�T{0.�E�~ ����2ôy=����D^'V`����.C)р���Yy�ƴ��H�T�H��-:=�nɌ�n]a/�X$B'~K��d��@N�cϪP�_���z����#�߁C,�XϷ����zneIFb�1����7�����}#��I ��i�'�*��U��!a���u��f������ij��mhZ���7��yI��dx�&."t$�H�H�� Բ�9�m�7�,�k�TL
]!��)�F:R
Y�2�9�B�/�����+�u���Aqyy_$�:t�#��_�+���ő��r�LUm������L�	��p����Svpȟ=�SH!b�GD*�[�|#���ض/����\Xx淳Cw�ϿYƃ��u߳�����W\tp�))�5�>���;m�-�W��6�zC���y�_����0����N�Vs�>c����AFH�!��9��Cy�x�������ۢ�WT׋��@�Z���h�vaF�W�?Zo�ݮ~�Yj��.��8���"7]c_�k��V�=!�>!�o@<j�9�آ�1F#���c�x�����8�f�8�ư7�GQ�G����� ��Tr��q����x/F�8t��Vy���*��k�;Nz����w�p��\bfcM�Sko�U��n�V7����J�jVv�pt�?�)ָD���n�\�o\/-���:+j�N-��J5��w)�:��L�W�-���I�,:��k�e�Qi��c�6�K`
�΅�b/g����UA���Qwy����C�d�^i��~-L�t�nX�H�T>��3~p�.�_b�mŸ@"d��п�Nwx$���5�����ǃQIP�������=�of{f���@a��RR���b��c#�\� � Qj�X�	Lt��o�LI��!�N�ZTy�]�s#�'zpQ��'����Ᏹ�[v������[�ܟ����?T��l5Z���'|��Ϯ��ȴGH<�߫W�E&&�L��ftv�i��*�F`:QC?�X��i�Iۯ���J� [jZ��y����VUw��� l�r���8�c��͆6�<�8"tы������̋�:���ҒB��쾔��1��쯟�|#~_�O�����8zGB��~u ���,��N�<oH��fk�|j�3��a{��ß|xu2�� �U��.���[�
���J�8�~�|�C?c����z],&:��_���?Egyi�շ�HS�c�QclW��y���4��Ђ�O�s�Ǐ�_�ҫ � ����`��	]�#�+�*�h��Oc�V-������ m1���5��ZӦ�<,��m`��r}t4�/<.�W��õBN���T��T�����d���:���F�蟧�'OHl1*QH����\h�Oa��U�����Bv&6���Q���q���(�2���@}���Ϩ��w�ͫ���x�끫��:��8Z��������Iw�/A鍺���,��X�L-�!J7A�t��p����1�1���E!ť��,�a�M����h�� aJcJB�Ll:u���5���Z���@̖�9�A�Z��Vq6>\�ff�v8St%]A��}X�k��78$�2�Q`*H� �n#&X�̹����O:��&���,��Qeyb(��ě��N�ھy'w��Fd�J�HOYy���_]���`O__�7�7���?�ؔcV��~'���6]$Wգ/+1#���Y���N�YII6�bΎT��������caa�����T�j�|VU���{��>��e��5�ڧ��}6�##uV 41{�0abW��������� �rE�()ޱ���1��{�����T�������v둈����@���rE�#�m��Λ�pm�qsjb�p����̡�`gb@P�DA� ���*k��E���vo�	=���Z_������"4m����Y�:&��i��|�m�%}�*�a�$�;��_1��ly����)���5Asȣ���臒�(	��e=��D��'@{@���N��m�A�O�]g2��[�T�m�`'�Ev^۶o�D�M��l<��Mf�ps+\��T�u��ؖ팊�rlD�^�;�"H�:�#ۈI�3F��)���rJ@�O+Z{D�������O;|��y������/zM(��֯�0��$(V�7}��h�ЫW̦���D���>���̪��Z7qW���H�Z�(ԁ�MN���㡡�X3K70�݇��������
�t͇���r-Dy�'FH�1��Șa;�[F
��ó�{5�xM/�"��:��a�tv��r�]�-
�#�q-#|��
��F�Β�\���*j7�=r�G�$!E��C�i��Lp�Ӡ�	h�[s�+ ���֢Lh�8Q��A���(G���Ä�G��R��,$;����3v|V{#_Y0�t;�-ꟃj�=��V������Տ�>��(��$1����!M��2r���i��MC>���\�Ș�<}R�-)�˶�P_�Z��	&�^,n���>��H7�I�p����:�j�Ս��������%�;�H
�̱GCJ�\M����1�����YQr!�߽MyY|�{��)�0���� ������C̱-'�JH��B�"׷e�v�FPL����(}�:%A�R"�_n���5T7���	�{�J�VH`��ǎ�`�.YNg�Hlo�j�)�b��5��w����@�w���S( ��kA�Ί�Ts����x��8�P��v찵l�� ����gO�I_ǈg�:(�Y �[���������`lO��<.3��76��9D�5���Y�����V=���_�|��n+v�.���Ș�~)U����g�5o�J}�"%ƻ�z%#��?Q�D�6���8 �U߇l���(��_H_�sW4��vfr �bE����2��Y�0:�=j|�R:�'sPs������nL����"�G6%�_U���@	!��3�M.-�;|?�����.�w+?I��N�*|�j:�q�0�2}W6�>�x��@vGvf~Rh��Q�����,1��`!b,[ws�R�W���w_vW4�r8��'���|��HUZ?�q��G8���������C|$"Bh�g�˓�Ƨ�eN_.�<�Ľ�%�#�t�^���]�c!fh�B��-d�~g�|�m�!� F����jϖ�"���~���Q
��[F��l��}����;��ng�ʐ��x!�6��s��(���@@�{dz�F�D�Xp8�CU�F��kd4_����9����U�ݓ���U٬�>���ɏf���k��o���%`����/�!���G�b�p�m�+#���{����!�8I��-ɤ�=�&sL2$5&*;��2�rdf9@��s
��Lo"P~W�J99�Q%�x:�s�O^��_ڳ���9|9��D����_��<�6�9D�u}�����*��	��vMpH�ϵ��J�b��m���7H��9�
���|��;eF�.��=c-�z�=�~\��a�E=��5�6p�,�ujz��X9dEl@�	֪mE�bj(ƶn��d��T��Lw?���	�j��/�A��@�[s������8|��?�K=�0��!+P�c�#�?Q���7�}�G��e|&_�\.k�ި'�Q41�tnmi�%�X�׺ :>�~g:ml�/;C��mD1M�`��O7��l����
f�^(q�2�~=��8�-3�;��d}V\П����t��Y)~ƿ;�4��~Mm����d��Ζ ������($2�w��{s��XMt���\������$pV�d��?d��0�n�+��������h~��dw�L�\j���2��6k�����J^Ȣ�g���Am����9���ȁ0C ��5�AYmA��Ω��ʎ����6�\3�� ��b���%�.���\�mG�R��)ύ ����S���j��zY�����jY�:����Wh�K�j��H�fw�í�>�3��.�¢�ĩ ��lJ�F��P(�h�cP��`R���"��(Ivh]�N�vs�D�9�6�8׽�t��e��(1�M��
-`2��*�kNSh;���(�#E��nm��`1�p�ЏͫW(�`Hv�6��:? �HT[� ��e��b��)��i[���4q��-6B��)�˖�j�+PZ^�����2C�-���̘���=�>���Ft�����k�6�`d��sb׬�Aa/�Z�2�K����oKO�\�al��f���	���2�9�8�bЄ��v�1����I�� �W^ߥL2~Mۋ��}�GgI���bI♖��-3�n����n�gffd�[[r�gH-�>.o��uR㻙Xm̆n�籓+��V�:�I\��^�Իo-S����>I}�� �N�z�|����?�QZ���ME�]Z�o>�8�T�AF8R�d_ɜ]X����Ĕ�(~#B�P�5�l�`���\B$�sx��M@���_�ְ�w�S��Yg0U!����*������3���w8	��66�a�~�y�"AH���O�kPz��#u�a��3:{��/�=��}���hQ�u�P����yQ� O�;��p�n���n�L�'oi#{�o�ĭ��`�m'���MD�
纟P �{��MKӞA��6܌�0�_�d����4�~'E��j�����?��:�%C͊��ј�1��߶�*:���N��ɀ��nͣm뙨���9�I�	��8��$8��}^��u����@��,F���M��HĬ�`Ez�D�s���W|;E���+3(�bN@ �%N/tB��L�W֍��U��}����ַP�w��0��$�c�GW��n"(��AĬ��㸰>M:��Y"'��>���Fn�"��e��>�X�?�P̓�����J�V�����Y�\A�'�˝���N��/�1
:���\Є�~�����B��sZ퇿��<_�e�i	
�WT�{I�9�>��,�l��p��yB�>6����{)L��T��$�2��q�ֱ�;'�l�;��u3��e��5<�øl?�[_���
��v!�h��ѡ�^RU��a.fT�r��L��w>/�q`��DL8v�Kx��/
���� ��|����r�߄�)΢[��4p�ɥ�{|���%)��?j��~�]��K�^ƕP;�r�5t��3[WT� ���-���b���łd�ρV`k���K�L\ǿ9� Uk�Jɘ�"����w�_�r��Z���_��"���}�����A�w_@A�n�c/^5J��5��(�(����������Cu�w8"wx=�-��ۜ�ؑ��T;B��_8��a��&�Y؈�6c��UGM�/|��M�\��<��a"ɒ TcÝ݆As���l$��]_:���)�R.&$e7�V��O�-I#�������?�9OΫy��BV_g���$O;
�k��|Ujr�)"�OY����T� �3>�v_��Jky�^w�ܯ�d���t244|��Jv(7����X�/n��ao���%�
�/=�U`�&a� ��EN���Z3�L�����V�f�I�RM_�{����ĕ2��\�g{%In<K�[�T����u�w��ԍj�ܫ��f�k�b̯��s�'d�]ɔ~��zb����9� �JI!1�5{d�Ϋ;��L�Xq6779������g<e��8�8�-��|��UX��٬�i7��w��n��j�}|�~�\��MD�n����K2�>�2��^h�/��o���U���:�� �a���ѿM����	�-{���Q�;��Sm��	�,�2570��5�t4�Z����e�$��Y%��(~Ta�U��l�Y�t-�+$���&�8����:h!���^����R��^�֝��ļ����[2�[��z-x�ˎ���3����
��ZΌ.���I�lT(���?�-�a4{� "�_:�C�Hrn����:�����cƎLgv�~�21G��(�"�Mt�ԋ�TI�ʑkK������໎R)Pga�9�?K���n1��Qb�Q����p̯e/W�r�oq�Mrd0b�:P4�6�6Y�y;mdd��u����@�⋮;�M�׋���Y�EI ����wz�� ��̂��b��759���%���+�%0E���y+;�Lb�_�h�:�'n�YԐ3����8��l�ػ��i����,M�Y��ʼu	U�[����޴ �z��˱�qw �O��$˘%1��U�=Z���KyIs\���a�AT���q�K�U����O�����4E�@�GԆ�W7Y�Z�v�~�E��ь(�t ���\-v�h������?��oOX�� 2}d$+��	&^��S�
z���W%��TI6�ݹ�Ʈ��B��]4{��ۚ�������M_�u38��Q����^�X�NJ��_ĝǪrCm�����Xꠧ}'���
�����MnN����5�@�к�S.�1�`H��*B�����q�V��PR�p��NY�"Y�����%���p�"pG�ر�"����,o�$��|vz�?/��b�����S���-Be�4�}��C�l0�^\�O�˝�|(~:�<{�8�w��E�SQWJ��i��e����#�F����e�vg8S{H�L���垹�y�o[��גn���>X��_e�m�ǉ�E��+�e8�,�w�e���D����9�N�%���M�
�Xg��tG\&�����:���S���ZwJ��`V5������`���(O	|�SV>�n�Fuj����l�t+���gt���;#O���6���I)�Q��*=L��7Yt�L���������E���y%��?�;o�9!�N����ּMvL^�S����pӪ��7&XMD�G�0��#����7�J$����}5�^O+�V��R&�b���m,��\+�����(gV�<ɗ�q�O�h~[�?2���z�/t1�)��AeX�U=��q"7v�b�L��ܱk����}6ӷ�Ӧ�dP�s�C���J�%�xv�_��i_R��Պ�x� 4��������9O�rz�?YLa��F������힧[1=(wӇ̹�[��q�Xn�_���)���gq�E��,<�����zP[x�_���(~��#u�����K���?,��������o���鵓��rp;���di�6�uߖ�,��i��'z�_G!J�&Z�&� yO�c �-��C����O�����z���@�jd`0��f�'���&ЕK��L� �M!-�
Ǻ8x��б�lW�ۦ|���$}����`8>�Vv[/������o�a�)�j��ʐk�p��ݷ���UYYu٬�mi�s�!�i
I����NŒ3m�fn8����Lj�r���?�0��=�����0G�����v`&΅�.�~���g�"�n��M�`����WY�.\�I�ę�p�� e��v���վ�/iLQ_M����d�������b��%��U��oD���(�e�1�����oL���9��f�\�FV�`�pJa8�[�R��-��������!|"K]��*''��݈�R�a��STQiN|������p.���]q5�|�¶bv�Gn}�t��������z�f^����ǰ3�.K�H�g-���M
�'*e�*I�̃�����X����Ј*�(1�7~̲�*�0��;}H4fe�z��+۞`u�������z��2�d�b���}��b�;�Y�Ԑ��������vr6��%Ec�j�ülb�vGC����Ǫ�~G����ᇫ��m�i4�H�����&D�)w���e
�!"�H�Kϲ��%p�8��A��Wv�C	GC�w;�b��r'�h���h;�DزÎb)��Oϼ���:��K��<�������;m:�,A_�I�9���J"���}!�I�i��\c�a��G�eM`׹\��F�J<�4�c�O<����`B)g���.m�T)��� U��L����R(����a=���H��"��`�}`t�`a`�)<�F�}A��b��Q�dU�̳v�e��;urXڢ��9�ja�[���i냀�f�ՊLK �T�.EH��0�_��mg��M��Os����G`[�щ�%���@�A2�y�����M	zD�Ik?3$��vK�X�+ևx�J�o�,4�M�Al�y˙>�᧛M�t��T<E�C��tV�yl�gx�/4��(�� Dc�`"o������x�]�$n��Y�'\��ci�w).�,Q������m�4����H���UZ�1�gZS�'�L\�w��H:</���� �=�_h�R��ZJ�$���e�tM�y�b���{�"���k�M�@�_�t��,�S��oרC0��J;��H*��6���A�UW�<>��Xl��U��t�_ʐ������/�&��U��x4�Jo���L�OҀLl�E8u�	]y��v��"����O��Ih!h���R������!=ɫ���.T�����=K�
����E�!p�>��aY
��V͡����1�P����4?��� i�UB�lZ��8l<Y��Qt?!�^�<1���	}/b��r���M2�m*�k���F�X����-0j+d1"�ܴ���F"�k�;,�b��'�dZ��f�V��0T�Q�MD��JA#�#�&������m�wg�ղ7�8G�z������n��� &-Pd�^$+�c���q�W����1z���ҭ�Q/��.�?�`� B�G-��:���D7�*Y���1��RJ��V����ooS���?��$���o@�F���;����˽����������"�G6�w�p��Vվ�Z���HT��¯Y��iY0�%PBŁ��J��E�Fh�Y�T��D�����9��ߺ�n�z-�J��P��`�5��*I�i�<����A ���������eN=�%I��'��n�vi��Oլ�7�/M"l,��˶�5U��cʌi �ϗ�������K��ԇnQ�oB�LD�Cc(�%���i�'��L�A
���a=A�^A�z%W	�{\b����-��)�F��튫�y�y�ؤ�3�W
_�ϐ�˧e��3����K~}{�̗��F�6�Dr)z]�ێ���>�@`�V����I��E�
����[�/��Q��Nhq>s���c@L���[��e�WM��&�K5�,��5�8:f����L�Ze��D1H�Đ�VS��.oYh���m7a"츭;����-��2ޓ�Q ���hׯEgT�O4=�){C<���a	8/�$XTm������R��{��oU*=�w�~��-|��E�p/�1�%dE�~j�}�"X����@L���Z֒��$�)�����w�hT^��.a��:޾+�|3�\}E��J{zߕbnYe�����%����u�d�zY���n7>�a��M��u9،bs��������qe_�ؗ�6ܝ{�bc�X��y���,Q��5����~�*{j��+.�y:P�R�~�����4%�Xc*c���[�?�Fݛd��g�!]"���*
�y^�yDab��?&2ꆁ@ ~���6Y��%SŔ���Zj�j먗:��^k�LX���ΌFd&��(���"ȑ�&4�N�V//wn�X�6��"����p�2җ泽t2�F��D�-�N�R`y�h��C���&��B��J��\�p�a
Г�qJ']"�@Q?#Fܞ�y!ń9�#�ȣ�ܯr�g�`"���2b�6e�N�}eK��sU��*�HC�{\[`JN~�S�[����wR�2�e�I7�&���N�ֻr4�9�|~5��pꕼ���Ld��e����e=�X>ۤ�e�D�~�ڒש�3�>u�Y�iA�x���Ț��Pņ!�f������>��+�-�<-���~�C!�3ud�zLM-E�&��&m,a&�?~���ǭ2�K���sjx�P�Ƭ4�7l_�5#ܽ��}����`�xI@�7$1N=21w'���ik8�a?:��o��)t-s�M��D�F�x��Y�9U�ґ�c�G��*�]n���f����N=܀=�ݡׯut;B��*�:|4a�r�Jv���m�z��d���}M�)A|V��%�ޏ�.dD��(�$G{��C�0�����@c�ckfCm���j�,�q�ؕ��ODW������{�xyʱ��r�t�mVC�Y[[�>�["�����e�rDI�Lx>h�f)b$�
�䄸��P�P	H�Д춵-��JC�@���H��~C�Q�K�2��Y�N�� $�����t$NC�b��i������\����s���N����!4��\����]��K�b��C���;jK�9��e�0aYz٫�/b\
2�D����ܦ�V�	T5J{�d�����"�L{J� E��&�(��m
�I��H��ؑ��_K��5_,s7/���M�*i���-M��n��p�(�F��0f�sM��^���W`	���ܵ(��!f���\̜y}��Y���������.�M���H�y��Z��r���P�3^������×�c���|�U!$��DԄ�]C�����k�Q�T ![��܃H06����5m�v�?��?��4:��{ro''CĨ���_
� !�@�!h���D�*�b=��}���:���v�?��Aod����1�*���p�t�W��6��W�B}���]�Ug�#�@�X$�n{�B����'�����k��Q��L>hkJ��Ǜ]��eљ�.���?�ޗ�ds�:���,�V��|�cǻ@�0ٖjT��&�L��ɆQ5[������ F	8�:޲��~�"Ĳ�HEnFu7��%&�I� L�@�(M:��S����W#��A�h�W�b���M�$D��sM�["[i6f{�I�ZkLo���H}��`^�Ĳ<�#�M�h�b:Ҷ�WH+c湕@�L�Dn�K�m�٥�����|(����	=A�Ġؿ��_�k���DX��`�p��9��[S1�7�Ǳ�:֛�^�.�|Tu��센v	d���~��� �|�+�_|h0ڹM\t�!��Fex"����5HO�(�~;1`��M¢�A8��L\�y�����>)���yg�3Te�Cu���nЅ����ں{n���#�Թ��q��Î��h�=�>Ky�X&�h�W����cIb�ƻ�J� ��"���`8��m�(i.0A(�@j��������vͺ/�+8�0�$���a�M���3Qڪ��a��t�/1�i];W�iVy�jS�&����E1��*�NU�2����.�����|�E��,%$�6����X�^�G@L��sU����ep>�T��+ڊ��/�O����!f�J�Q�g��c�W�UVp��s�N�ׁ�|�(}��`q�����C,^�د�<ܫy��?�t}��7W㟲~^֢���{������>�8����DLR�*�ΟTs|���,{�w�Ͷ�TZ��]��@���q���F�!��h��^/��߽��k�c�$����[GfNS%��,��_���b�Zj�т�4�$�Q�����j��>��?��}͈�lDk��)����|~���0�uob:���.�������[���K��� l:���v=��mۃlN��2Z�k�>����d�v:��c��GU�t��j��]c��	�-7B�M7����?C���pl"�yK��QkM��jO�F�G� �'1b�=�I�8A(a	��O��to����yxZ��5n�o�h�����d��)P��+���|mu?<�Q]XJ��#��b��$�V!U%1k��	�ݻ��lL�`�3?�,ME=>>B����;�#��.����U?qG���c��/��������������Z.kr�*!��$WE�X�[��ۉ���qm�oa��n��[���']�I�AYϻTй��WR_�*	Whuw[�#`;�`:��Ѹ�'p��Lu�9����;&�
�x���F݈�����J����$9��]�$����Z�A^n�il�0~��0s�G5�i�ʻ�y�ϯw�k8�F &��[��n<��M9�s���cQ��(\��0-ڣ.o�9q��(7mh��,0,�!�KաM%�0�-���$���j�Xv�܋S֪��w�z]VQw�9�ʧ�U�p��O�U<]٘WR�w�4ef�'���4Zpo���J�?,c�]�gX��{��>��}#��T��7���
�LV B��%0V��?�j3!>�D���a�k_c�eHs?v�g�O�&��7�$z)�B;��T�������~����I��k��J�Iݎn ��xa���c`F������m+�A��|%\v�d��5F+R���w<���t�"���\�{>@]Җ�!p�\ť�
#oC@��f���3p��B��L�L��d��i'�l�J����ٝ�d�X��G��H��$PMr�69��,1`���Q  ��������oO��9�p��8z$�^l�:�}*K*��{�߷��?��6��ǿ2��:�~56�D�8t��[�N�b���a�2�9@��
��H�@4V�T���7����^�W$�̢t�&�����_�
1\���1��3�xt�Q?�D�W���r���p&(FO..&��9�z)�!>��0F�}uɺ?�?�o*E_�{���1;ܫq��cG,��,���R��`�XII9���a[���-泤eL�K$)$Yl�v�&�PR���*7G��W��F%`{��whr6T��q�0��T������e�+/�~M�D�Ғ�ko�eTb(�RM�ț䟿N��F�]2WK�d��]��3`l_{E�r	y�C�;L�p�����m��FT� -!�7�"�n�_��ַ�h�E^ΨX/|������2��������Q"豞��%:
�)��S�Q9����<�~�*Z���M�	6�=��_B�����͝�ۉ�4�/�Ҭ3WR������7�@��VE��?@��ܖKq��5Y�t�:�<	��h�F�0���&��?��XG���GT~��w���Y����w�?�~z��l�_M����ۏ{�O��^lbVBt_�;a����/�B]~�HG�>�	w7`"���ϭ:��[���j׭�+���׫���紋����3�4�������<���*�,`��_j�z�6m�u�,�q����
x���P�+m��r���<���*M`:���f��D���e!]/>h\���I��/vO��Y�������BvK)؎��Y�΂�C��M�]jgf^����W+:fM.Ic����p�a�_�[��8�}��  ��j#����7� I�[�*I����L"⣣#�#fU&��^dMB���L�*>�L��L��ZX)��N��|hjĎ����E�4?�C��.TO���ȘCm�-F�0Ϋ�)��]�C�6y<g>ĠPϷ�{l�MW��㠶2��w�$�Ƥ_�+�88��V4�V#Z�2��TʢT��U꒤6��a��7�8�� ���ˉ_5�$�!:=Zv�_w�T]KΉ���_	Ձ�hj�k	X��K.z�T<���;Ey��Ϭ�귍/o�ȡV��0���^���\V�f�krg�b��t���aR�����D��ڡf�.z����@���j*d�Y�h�@1QnBvs���HO�����s�+F~�Јj`����8�L?����@Щ +����#��+�dP�x���i��B[��IB��8�{���纞"�/G�ɵo��K>�1�i���P8�N����eͷ|�T���'�Ef�f�֎��|�7A ��7�����t�$���x�"U�:�#�������~��μ����&���}Q��g��;��*���$�VVP�aݝ��xz��<w>��ﶌ��Y���,����b�jCz���+���+B�q�tNU� ��z����]Ǧ�6��`F��d;��������xٗs���}�*i��W󥹸N���Fd2�f�D�F�B(��O{w/���{�!�vb��k �[�zW8�7��?b���u=,?�D=�8�V�K��l�K��}�] 9P�PIZ�8{h�y%F����^�UcZ��E�����瀚���i<�|܋3k�h��C͙>8Ѓ���PZh>�B:iu{�g�% ӈ�#�I�4�_}�����3���8��ҵ��ǫ(��E>a7Kd��N��i>��cX�r���}X�(Os�\��{���lH�zA�	;Z��L�šE_＝�Ma�;����n�ʦvx��o�űD�
w�i�Ǟ`ԁ�vw����}�JЁ�P�ջ�S�$����:��S��̪�����[ ����5���{qkq)�Pܡ�kJpww)Z�%-��ݝ�,����{�o�f�@&���=g�yvՇ��ً�ӡ�A>:.��\i-ч�������6�~�>�|#��B�u�{���e��u��~a[�������X�Kpmwi�P@�<�_=5]����T���%�Z%�h'a��+Sk{,�t�>��z21�q��5]D���B�/&v����g�D�|U7\R,�S������|���';��
�R"�{8 �z��4���z�~j��B�^�-ϊ�f����r�g+� :�NL鱸�G��h�q)ܳ���k,��m�C󂧺������mҏ�P�`Ņ�m @-�q�T;@k��P��B����u�O� ��/�#���%@ɻ:ߖ]+Y�b @��£�
Tc��Ƹ%́�q�r7�h?����e�:�dP�7ֵ�u���{��Ġ����:��OҤO�$}d���-GF��]�u���R@�W�����wZ��PB�3F�m�?$&��^�"=��* ��?��!�ġ� /�,T����:���&���:Ǜ���]� {Lç���@_�a���P[&�쨳IQ!iȸ��?=!��ݪ�eJ�n4����?J 'YY����_<Yxb�bvSu3��MW!�:�]�W��X�[VP�E=\��f\.(n�o�+iMdy��F����X(�a+ÑU_x˔oR�f2�EAj�%�<UH�Ǔ_!o��$;�����Zi~0����'� p��%0�X�'-2jo�_�&M~4�#ʢK�o���L҇#y׻�Kx1u-Ͻ��I��1�^n��mt���6�solQ^!���WS_+n$���T���|%6�)'�f�:b.!�q�2�ٰ/;>;��Z3S�~��3a���M�b�����xLV���#%���ZD\O6mmm�+;=�N͞�*�L�e��K�oc�a�Q&�]���n�����N�L#|����p��beh���)�7I봅��g�;^��QB�K�a=N��}�}c��n����!5[�>YMw$�@T)�~M��Ǔ��t{W%��&5<o\V�;?Op��˱lFC_^V����bk���)�o�Yi��������a�ҭ[���6�y]��VL@d~��4'�h��\���4 ˮ������f��k��*� (rI���ș�H[?4�%�k�.b�q��9@�,�$$Db�Ͷ����S���c���?���x�F�B�4hs��[��b��c��fA<lZe�]D�s� N%*����\��a���3��-2�O&x����F�bj��XbA�{�ի������G�c�}�O��(�J�F*��=�������^�q��毋����:j4�m�߼�/=����w�/1�w�
��7�J�`[��b�8݊���\v<pW1G�\�E��o�`�v�eA_����L[�h�8{�W�p��?�pt���d���@�3�'@a
�5���<��	1d6.F�&ԨMYt|��ס�5y��6��<�Kͣ������+mF��&$֖s�~�?Tl�u�͘ޅ�U��dj�ߨQ��v�T�{վ��;�`J[�;!3"nB@� ����E��f��U��G�AA!�j/�Ȍ�f�5-�g�n�"}Cң��7-�R�/?(��/UfgcUt��,V��}���?h��~y�����&�
�qC�2�4�9�~t&5.߹1�q�%ϨLY]�����$��p!�wc��Ǉ��+���U#pA���Ô{�2g�0(?U=����ވ��4x�[�t��<�s����v�,حLH�s<��vv���;�GM1�晭��	���#�0H_�Lj�ޖ}T��`S[�	�\���~�6���_8������R��	Q��f�Z��Q�/d��1����7�}�-�\/K���$
x�T�=���i��ϧ;�Y�y�e��򰆽f�W
M�q��;�_V?�'���q|S�F=9����X򾇺ެ�Pzi]����:)��~�_3�#�q�fX�5����� �U�k�����*�N͂�d�H�#����H���K��&�I�����+��W9N�W�
��ڻ$m��6
T�����t_�K�V;m˔��3OV�?�#�y��-	җ�c�-q>���8%[�5����հ5�񦕷���Ŧ�@���[�?0�呴T	���)�d[�E����NE��Yz9�_k(���m�^�*�@$�҃����s*K�ʁ��³M+K�Ll�R8�3�W�~��}�X�G��k|C��mAq��5���@)4�[L��U&�z��#F��aJ=ת�L��병O	:�[�8]�m��Ǹ��f;����ϪY�nN����ݵ������-)�H���������-;,2�\�w1�YJGG'7B�,g�[�_�{�D��YT�#���<飂��H�Wu�N������z�`kRO^(�`g�#��6� ��\o�]�ջ-
�k(Ǹ��=�-1H���\G~��*����+C�{�W3m
��#�\N��C��t�[�U�1<)$3�f����\��y%Ve�絫�N�H���OW�J�6��izf�x��V;o�/� ����|nl�7_+^׬��n����)�ՃW��8򥏂�ҍiE0��`#	�غ�^k��a7���	{��=n"�����nK/m0����k�^�!q��[7�)J�& /F����TF�ղ��p#n1_�Ga���h�2̃]�b�\)ac�m�Śh�Z����H�@���G�beת:��Շ�@U�)X�x�YUF*����Eh��B밶=���=�(�N�E�������L-!Td
c�5V͞Yg�3��@�|Ar����o�7����uy�����R(��^$1��K����~����˥�:R��EUv�ǉ!3Z�����9}��7�>�Z�FR��s��s�C)#���~�m闆{]Eq;�A1���z�;n�Q���b2���A�PV+���/�͏N.�Ə�o4�OJ0Q{�W�	��/6��]�5�C�t����,V�2�x88�1B��0}��Y���z���P;������Kp�w�D�_v0g<���})��Gv`�YvXT�HL����u�#��$'"؊K���C������=� s��?�;U��Vّ�|���m�����{y�~<�k�S��b�*��f��-`
Y!\�gq!������F���BTID��Q\3j�;���Ⲫ>���߆0�7X풞[=�7ܴ��!�zRsF����_өw�V|��Y����Zʂ��D��Vg�N�yHM�g�ʡ�#޺czԪ���*tg��'�_)�pQ\C=��K� ;�zъB��j`D��R�^D:E7r�R-q��K�}a��ՋA��q��vV`�<3��ǩ ۷��I��G�����b�����q�17�]��a�p���qlVW��/ED�x�ڴC�p�sn���2���`85��g�p�6ᴏ4; ��[��C.�w�v�
��Y�QtQD�T6���@�2��Cy�@�e��$JGn���)~�ἕ�=���p㸭�Iq����M1��E��CGۄ����M�g���蝡\ ��5"�}i<�R�9��[�nHĂH}���1���{���FiYe��a�M�Nf�CꎓC#&b��z�&ܡ��šZ�'|I��6����L\�Yd>L@|v���x+��xN��Ɩ��}�kOW�h��d�> �׿�ϸ<�4��8�=�'�n�|���	$`/��z*v��m���#��O.��a�E$$R�v(X�#i~tz��Z_�8pF�I�e��D�N�#G��{9�Nת�\s�&߄S�<��r�R�����}�`Z<�nò�2]���#��|>԰;Z�哮�T�R!~ʭ�'��x�Yԧ?2Ɋ��8^o`(�,hz����ƾ��w�NsF���,�7q៖cS�Y{���� :qoٟ�4<���8�D>Б�U�Q�����H��:g^R������"����)�3�r�wԙ�k�/��0�����0̮���g#팱�-�I�#�A��E-�C��xp�F|z�r�IBv�t� n'-���pc��&knYӊ-���)�4)�
7KM ��,nE�]�|���@(2�&��hH��p��x�O,��;�v3�}���|�e�G����Yr��?��n�}�br���C&b����\�����\H�	Uz���ӿa{5X�T�1�玮<��N!��\�ђ���P�;d`��G�J�Kj{�c6N=��C��`�,g�����B����[�B�f]�ն1�̑�z���˶&2��Q��!K�������⛿$�\�0������8��Ń����P{���I<��|R�"��R�� �^�>��
��qgnT��a������[Q���l>�6�� }��u{�.Ζ��m76����kvJ�;(�QWzg8� �""�F=���云���^ZQ~"K�/��	���d@���
�QGX_^e�`#1�BL5��_�ho��M��d6k�z�J�	&��N�o��eƭ���$���i�'�t캊,�D[�� �V�:*�T)J��%�uR����sP��j��-d\���t涞 �2;ӏ�������9�����u�Vv�^� ��}��R��Ŷ�����"�|��g�;V�9�ȧ?�+�N�r(agL�ǘ�A�+cO�\�R�h�����6Em�������c�K ��Γ�7�LKY(E��z�9�%�]~��G��j�w۫X���k嵺xc\\U���ى�����z��P�c��)b2�N�Z�zN�-u2��A�m�|���Mn�݈[��1����r� ������$���MFOꒄI���U��+NS�,0��N�ER�s<��4�5���G�)__�E�	C�>4(��e�!(�_�O�7�DG��$��>���|$4.�q�=�^�w�Wl��j�$���	�9�?xUk)�8�t���0Z��BwN����'�P�GOuc#vvۅB�M2���I���D�1����%qv�-$�&��ӝ�9�?�I�N{n�U��3T���ǈ?�&>^�d�En&�Ϗ�c�Fd	#k���덴Y�w.��A_m5C?�%@8U(ϐ�c%%:���ٰr<���9{�ЪSF���)6���<C�PΫ59�3��w�b�f",8�	�k�ǉ_�
#k�CaӤ�c�&�GP�{C%����������ڔ���쉚�ĦgR
�̽���h����P�7��a�,X��/f��'w(,�Q�_�
B�	����v���MY�j䘙�_�``��N$�Ig�2m�ǖ�@�B�)��|z%K}��70�?���H����9P^��zI��І#����{�#v���vE+���R�8z��sxff,\�dco��z9򧐷k7�&������Z�N�JWK���?�y����4���8�HC琚FԫD|3el����d`Ѫ��1���tw������R�����l��*�s��]L��� �'c�� ��y|M�%��B�Zߢ,w��%'�à\��߶%}�O*7H�J^_~� �@�x�^eɗB�	j ���A������{�{yn��L,N�X����F�{M�%$�k%\��kx��9��<[�>��5�8OW�,��k�cyܥ�տ�*i�����w�۷Ǟ���pO��G��DR6ז�~�����Jl����5t�"h�����=g�1�Ỳ��$�.�����WYMm��]�n{��_�ǅR��?��,Q_GbL��JO����]�+n���V]�L��r_����b�ŕ<f� ,!�dǏ<t'uV���ڡo1�ߕ8��ё���L����Żk'^�*����m�߾*D�c�3�
x1y8L�M��MH �E�=�l)Q�ż�Q��R�b�vL��(Y�d����7�T#֒:�h����9�8�[.*98ir,am
��4U)r�)1`�"HL�u���[k�K���%���w����o������Ff���,���ʻ��{�Pu*�d/��g_�n��@ه[�;��,�gC��K��"��Y�U�vu9F�ʵ�~t�4/��K�B!z�_i5/T�(�������U�G���(<[hÙ|�fw����Fh<ϿGv�]u�����Q3F���cЊ�������P~j4w�:�;`k1� �	��'�WY������(��C��n��f��t+�3����J�0��(,��C�rSe���s��.NV�/�/tU�>�P����禱�~ݱ�"�� Z��s�;�۰�f�|s�]����"�i=�J��5��@+�h���%�Z���ۦ:��}hPА��w��K%rj��,��2�(vjLzό�޶Z�lv_1�}�g���Yf����yߔ�6�Wt���!y��0*p�DV��w<��-�;�C�y��!�=;��4�䭞���&j�g�smޗ�r�zA���ףծ�BV��y��}�+r�l�9�ס����&2	2��*�;J7|ОJ�^�题�)�Ņ�����f�75�D�S��J��#��i\��8<o��0vO�b��D��a95d*Mj���Q8���/	ur2pm���o���;����bZq�K�Oʕ2�v
�;�}z��;y��@D#����z('����s�|��`��IR��z�k�m*��lTb����c^�?���K5�G����Q#��M���k�,�Ctt�0����K_�vTX��y-~�n uT��(Oȓ%Cn���{`�w�|HU�O�>�>�������l�uޑ���R�!ڤ�
�p[�*̋a�y��0���I**q	����ݪ�B��>]��J�Y&�\?̯��8x��ޫ���jH�Jcǳ���S��w���\t�%��Xv���	ؤ�Zk���h�� ��n��B�y-�l��G�R��fUH.�+���J:,�=�2A3��Q�y�Dag��;�a#	f��B�kn9�[L�fܝHڮ��6�Rn\����=����^]N��ON�z�	(���R�֚�x��>���m�� j��р�_:�����|ܹw�zTw��`d��٥�[�[�}p��bo�r�Ţ
A�� �_����+�{%��K�%I�>��z�'��>��H��L��vİ��O܀Y�]�� �]���d�~���A��uEԹI5�8o
ư�d3���@���X7̡F��!�s��3��#��[�h��p@����O$�"�zK�Y$�N&�A�%�[@�Pl*����1j�*V��ݿ�ݘ�b;�����;O�[�]�h�J�k������7�AT�:4b�uX%���<�,:�r����_���u��Ц.���+�ѳ��lq�T/��=����ߌ�꬚y�rȲ^�+�@�kUm;1;�?��4�
�G=�/Ub���i�I\�7��� �mx�
�O>Li}�A7Y�֕���V�z��x��.��$1i@J��#�S#�!�Ϳ�J�=����̹iJ҉e$�SI��_Bޒ����Wc�M��-Y�������?� [N�.Eu��B���}����3�[vl�7�ߞ���q��/��foVJ��q�|Up/�'�& ��nO�����{���2RF������\g���C�uB�����M�3���>3�|/��O�A˃��������B�>!������l��YA/f6�{�3t�k}P�}��x�n�G�/Șo�~�%�@���叇#lw����]��|�'�]�ln����p6�����a�3���,���8-�t������!�"���@TQ����Ԩ���uL���9R\D
�(i�ǣ�ܟj���Co�5ҁ��!,��l��������:���m�$�����v�r�,��������V+�hu����5�a�WY��&=ۖ!\����3��`�f�jX�Ϳ��9��w��H�T0�'9��*u�JX�z�^�����<��eХ�٫�مg�A���&x�4K�A�Ӽ�I��N%ۿ/��ĆS� �i��l�9=��
��gT\$��,m�G>����Li�Ù���՜hL�O���V�E~l�1�}�� _�i�B!�/��M�Ԇ'
�4�3�x]��C�evڲgdY8/MኞNu���f;7��d�k,%Ql��	����ӐA��ܲ�ё��4
����p:jQ���\=߼�c�8�q�Z\��	�;v�f��؀=W*ms�"�Z~�s�Uםro��*���1aeC���X�� ��E���&��sl�o|.�D�ʌi�5���v0�7�ϻ,�����.^�XyG�i�g?Ix�]�5��R�\<�:��ԃ��Z!�
\"|a�6TB��>�u..����|�,bS��A%�Zc>~`�.�j!�p0En��_�j�����,�:�w�w}�M�S}�D"�8�g2�	f��0Mz�T�s����b ��䫅��'f�?��
ِ�O�S3�Gm7��W��ߩ�� �G�O���dn�2�́ATF�W��ZחwH6y@���L�FUp�$�?K�~W6p ����P\SM����v�՜x[:��L-��8�2PW[���D˼(3���S�:� �3�R�y�l�9����1�����l����Jw}�ne�mS��	b��0Ŝ��܀D�.��T��w��c�,R#ng�VI37=��Dzi�gtʦ�`��$(���D���Q����A��68��i��-���9*ĵ_�ݩ�	~.�D���<`��A<�Z�[ً����S�{g�&~�c�Me��w��Fv>� a��7�4@lIi\\ ���X�SV��Ͷ�zN٣���,�̄6@��=e<ZVW�YF:%�AT��9�i�(�g�z$Fa�*M�qP{�\�@�$�j#��ô�oN>��IO��sk~,T샴?P���Z��k`<S��Yo�G����b�S�Yئ6MZ+�0=7���J�GYĹ���]g�y�
X��Vվ�]�4��j����m�t3����01(��|�~��d> ş�0�dp�;�OU��17�ă_��`���(��~���kμ��Ac)E�y�x�.}G?s�:-SEQ�`�_������Vө��Z���te������̝=�͋���8�����]����W�u{�ƻV����G����%f����2l��}�#ΣVbv9�󵈋;.�l9���E������%9NگC,:T���7�d^�w���k�*ͺ�#�5�����>�oLd��c4�'�՟J��D��|�$��4����̌V���+�F�B�4��q{�o���g���5悃ˋǩA�	�Dq���aF����b-c�b��/ʿ�p��g<J�\őe�9�C,���Kf#�������׎��d�h���E���suIh�X��|�pUlqqr�@�Y�A5��ʡ���T��I��{b��lC�S��m���g���.�c
�J�\�85�f�����q�h�iz
����]���L�W��/ҽ�ĘUsjN3�	 �E�j��v��ǲ�ҩ�-z����|�11n1�g?22���T�?j0�&!���L�fF
��8:���F$Y��������t�����੠���C�ړ1J�?���7=���Ό�L���9�$�"J�}ת��QD���ʻ8X��+���n�TW�r���0����:Cݺ�������P6F�hr�DU}Ԏ��b��k�Y�Z�*۟�r/A����}�	��[���c-���
7p �%+�aE:Ψi�_�s�I�r-��
h|�=�B�r,WƏ]d:5�8�����w׾�y����7r�����:�\�-�0�)��$��K����j�����<�)�t��<����<��y�M��Z� ���$���?I:bĚ~����^����.[��'�sq��=#�o�r�V|UV�ڤl-k���G�V�_�f�D�q���j�+W�蠮z��l=!&��L��@�?Q?��C�9K�����s��L����Y����<�Ǩ�wF���\y�f�(M媂՚K�B��3@�(=K�Ҝ���S��w�R"���uY���Aa��8�8�����*�a�d@+q����%lR>�	��������� l@���3!�B.�]6�Ԯ��eI3R�p���ޒޭ���  �9�x\N�H��x=�)�Hn��o����lc��u45C,���&��~��cqXw�z�zQ7h%�
��w�@C�Xo����7�~�C)y���Zq�]0�k�	l���������zN���Z�''��4r�$�\V�C�6���'����t��N'?���Y�+���C�ٌy'@�(�`�]����n�����$+T�`/PG���c��u9ca�^[CCc�0^�σ��韽X#�>c$c�Ȑ.�r�{u��c���b���|�ujTqMmMnELe:�@��p����i(Ԑ�9-�t��>YG�IJ*y�� ����K��"�6�(���!�IJn$�o����|�e��o]��ܟU>Hh����#�o9����g����un�vs�	i���C�i]���d��]�r�,v��~`f������u����G��|���
?'��k�=��������)�bHTI�. _OC�6E����Z뫵���4���}�,P=b�e�=:b��y* ��8�n�Щ3���s����x����yl��4������7_I 	[�2�����:mv����o|rm�����w�
�������Lv�c����	J�o��w.�)�w�=�5���Kk� )B�}�g������3Dw����
_��D5�q�)X q��H�َ؎z�2a�Ҍ����?�'��Scm��
�i��`�V)���}�lfOc�&$�5��a?e�h��!L+��MĿ7J���׻��ݐ�G�L=��2b��_���8��(9e ��b���f��ׂC[��0�r������v�M�X?�t2$_�y�"� You����s�\4��\���榿��8�fe���"�(�W��<=������ml�io�zI�9E4�"�|�	{��M��Az��1}�1��5��mơl�jv>�}�K��#�q�N���])�6�����D�� ?�����������=���EG����]�VX�p���*#ti�C����ON�N�}�٪���t�؜�`m���:٤���1�N�LT��a݇�e��s�IO�>���aQ��pC�-�w݌��-VS[����~+x[R� P���lix�&ix֦ř�B%5�l������e��cG~����z	����w�+���R�?� &��@s;X�w�1���c�
:7k��t/Me��Y����{�t�RQ���4np#6��ȳj��QU��xޢʆ�[�oa�qE{���_�M�O�P.�u3i����'���}b{G����b��n���Q|91�^W���I�I�����ާ}Dë8�'Q�J���Rd%!!�$�t���+"�ݎ�&��f#c������LV�*C��9�X�O�9���3�!�w����l7�bGW��:�R���y`�)����Q�]��$?���5>
r�����M��TN/8��+�����N��-���l��a��X1p�e�^G2E�5���t��ިT翇�-dh�v�K]���A���{�iǚћ��ޜ�0��c���ۭ���^�~��9���W&sC�ӎ�X��j pl�k��� 4��AO/�i�&�y&@S���	��� �	8be-��w�'Lԃ���M�~���H߲W4r�l̍������:����{ai,݋-�m{#-D��V	=�2	�Bv���M�_����M[	sCA�T�D��a>��A��}}�yI>����γ�%���S҂�i��	�z	�X���ςM)N���G��>�g�=ۜ���^E�h�oj.8����>�2˒������E>.P�|Ssh']�}����1�u"8r�����ʬ4M�4痃lam�tV�;�[�9���6橡����<�9�0��{�lfe��;����<ԥ\�&a�/����8��Ⱦqg�'\1Ps��`��)Fl�0-��&��;�$АE;B��΅$B�TY���#L�hiM1v,w�v][�{ ���6�Ö�B6����BV�PʅK�ۼ��W�sBH�'|ָQ�u]?��e���P��o���MZM�c�Ӥ��W;��E�xg�WI����r������Ɋ��Q�Y���))N��M���	"YB4�hi=a���JJ����O*��~���t����z�)d;��X�s ap_�U�UwG9+8����2߰c4�opru��D5���E���"���	`��ky�"��<ݴ�&����+:����\��ؐ��g��)�X949�����ڼ�IF�mWw
����N?�4�M��v�b���t�N����_��֭��W(4�z-#@����}���Q�Pt[�%��zڃ�8%ϵ^f�h����&��|:	[v�G�F�}���XG&.lI�0�R\G�f�{�}2�_�߾}�Y�3b<$A�2�p��H8wXi�˄d�9���N�K�~,ϻ$�mw�Q���~h�ӣ���-���N
tƴ�_^��������?���^���U�y�r{2���=�a���r��qO8�|����� ���a����o�!����7�J���{ay�T���Š�||W����F����4r�2�)�{־����"姯��:+���!���~ E��-�-�7Yr�ʧ���F����%9�ϵ��Ɏl%�B�ٷVu�ƽ1]��T�$R�Ĉ��m;|�/o��>�4���T�	z�|��RXX(�#�i�ьF��t���B���"�k���`��۱��u!ҕƳ����FP,��?���ܫu���.���|��+eJӈ��&�A���v���,i>=�e������O���i�Em*�^�hMV!�%�4g>;�!�x�*s$�Fȓ��[ʁ�bq�K�������� �UQ~�a��\L�$����~лSM��)g�R�����y�H�BX
��3|%�!���x\P����(Y*Wr���#8�xУ�#GKvc,KvRH=�J����(���J7
/���v�'����M�p���Dyp�sI����V�gQT��H�¨���ԣ��y�[�/:�h����	o7ܾS
S׋��b-�t{fQJ�"��W]&%v=a�U�2�ý�e�,3)�C�i��A��]�0^6�M���*�]�E��������;ڽ6���]���r6v��{9���Xh@�>�5���Jb̕7 a���J?ͮ,�%ē{���Q%�x�!�x��?G��*����{�Y�^�ՖJ�XpBg��f���pa@�D��9��RB�KE�V/��D�!(tJ��nQ;��
s1 ����-�B��+��#�8�p��6�"F������aQ��7�#{i�R�G<�ixa��{T$Β��J��"��0쳔H���y�y-��E���!	f�?�9ԓ9�����3}���󯔍�G��P(����q,}�p�
I���9�n#�N�]TdO��_�z�v->z+�k̔�ofTl�da(�UƉ���Hwc6$T��g�R���t����T�����ow����ߦ�*,���\����{��!��r��p�^�,.
����R�bk��� @�WL���:��Ǹz�鐷�Q�:�����7&91~9l��v���Umm���M�~(�� I�V�-�#V��B��䥖<�'n� ����NA����m~�J�0B���p���`}zRUmq�M�s2~a��8rUT�r�/�c�T"���k�<�l�R�]���y=��23k�aYGo:ƾ�TT�s��Ė�Q�/H����iV3U�ᘘ�f���1nbbAo�A�� Gz������W[������#1�V�� �gٔu�e����I=����2fm��8
a5�4d�����6 mR)��_[�:4��<�qI:�o���Jlb��uk�k[��0�J��4%�����?@nM;u��x�%砩�M�p�.bu�q-GS�r��������D�g��i���f��^z5������3��O��\��yb���w_�;�Aٷ���ӓи��`T��A��}���G�$�&���u;ݿ:1Z��2�`�?$+��C�f�_�H��4�'�)��"2�b� 3��`:y��R���;p�Se��q~L��%qۆ���w�&L5�1'J��n�u?z��]RTV���7K��]z�Fg�IoyQM��'*���?����Rȏs��n��U:�>�x���*Y��ъr.��2��g/�Ύ"�Hl��e�Zp{��@!_��sP['kI���q"~�c�꽥;fLV���4Q	�S�.E�wq_՗��߀�R��qY���8z{p����kc�#��ԋ8�lF�d��Ǫ}�FW7�O��m����-$����7��U���I9(@=K�����܀�&�0n�����s��t޹'J�A`U���l$[��<^:��)2Ǐ���~�A,A遁��I��p⩈"��4[��F���g3M]>���H����sf��6.�%z0�`���y�'��"E�B|��� �����@���{�/�@59!u��_��)�C�y.y���zY�xO|e�����P��+��	E������Q��C���%ũGtU, 0w[^^^dd�?��Ӷ/�)�l/#L�".)iF��@�vۗ}Ƈ-M"U��p6��x�g�;���̻ھW���o�^�� ���e�T�8V���I<����vjy��,��~�e��ߤ�	��a	��6c�u~r�v��>��j���$Sm[��D�<�h:�hnwf�l����+u���k3q����a۝�r�E�8�� " ���+z#��y��}t��drP`���^ ��|���p�ij���a(����~
�s�f]$Zf»��R�a?Gbe�m������d9�mb�7:�`	1{�
���ge?�q��T�en�;6"����H��A�ڹ�E�a��O��6�6%-�Z�q���m�ʼ�����5h�8
�C!���6}�~~/�_�=^	�πږGo���cWBs��g�}x㚥bGw�p�{�kG�ϰ{����#%��&xiCG�QZR�o<�4p�z�߷�fPDs4}����\��p�}V���!�2��q&!������c�51a�{�^<��\P~)�;Z�\��T�;�7"��J$�����A'�uԚ���w��+������ ��T���Z�o��6k���V�m��a�.���Oe��*Gv(��m�;�NZ B{f�IL�M5
�K+���_CP��GYM/���Y���5�A�p��9�2���,C˕];H����sa��V;+��č5y�T�R2D<��9����Rֈ۳G{l�in�?��YYY`�J�(P�S<¾��������PFgE������p紉3���;gu%o�F��B� ѡ3�<�ٴ�f��iPم��]�#]���뱈.N��7L��uR�����?QH�͑g��faW0>��$M5N�����P��AQ�`��+��ΰ���s� ��]�}
������>�fFs+̮3��]�p&navz����|r��h��.��\����

�i��BLNګ�z�Zgf	ܰ��è�mѬ��6��&���rs{J�h�kT�9`��<3F��Y3��2����!��V`�;�T����2x��L��Q���f���ڴ�чn�!RN��w(K���`ܞ�%.�,�e���]�Ȥ֟i關q�_6��@��_���X�2���N��;�+f�S~Ȳ�E����g��؜<��sǐ�8�� �Q���i�Ii��	���)�U�4��(����-Va�7�yG���W����ĎS���<��Z�����j.��m<ߥX��O���d���.z0���չ��[���^~6��z	���Gm�s���V����6
.���Vd�@y�,\���g� 2�t�$�12��J��o�O_�7�4��\η�f!�6!�����c�6�u��^�Lgy�I3+(�	��P����-�Q��L
>�96�1K뼱AöEw2��L�\���t��A`��8�T0��PK�I������:�_bđ>�`�O�Wq�=Bhi�C����;i֨�"Lp�@Fn�q�P:��Z�����Uܬv���bw1�<��[�4��pFRLp�qd�G�y��ж�*��zH�ٺIn̚y3Q���i�֛�<ՏZ����p瀕�|j�B���1�z���8.��:n�Ȣ]߂yUX��ñ������l�u�[��61�j)����;�ST=����	;���w##sϬ,n.�/!���D3S�Ӎ�v��������$�4	�
��+bNG��D����+Z��a&�#�?2�.j�9��
5K���fA)�m��մ��b����O^�a�̈Ƨ�)����Ւ���أ\�͊�ݠ���L�}V/����R�����46�]i����%�;z ��(o��a�&\�И���hљPJ&�w^*<ĸ}�BRKKK!�����$���֗^7XY�rN���wY����Bحu�7 �!�w٠�t�K��.-Q���H3B�N�Qc�[��AD�0|�� ��F"�z-��£YL�5eE�É:�y8!|}iڻ����L�s�z�c�:Z���eAg擟v�޷u�����O_�v�}M)������w(P�X� ����
�X!�J��Z,�]��~���f��2�d��=��wם���`snڹ	�;�t�M���|G�pN�T<��U&QLY�Qn�2�9[�_v ���upበtC.���*��u����Ȗ̯X�B6��������V��\<v(�?|0�ܖ�r?emr�:����1��AR��8��ܩ���OVPo�Qg��~29��2�\!�l��	Pe�"�hn��у�ќ{q��稡;i�,�[�Y������+�� ���O����6z����Ӷ6�{�nٿ��K�gu�ӂ�?Q'~�N��3�"3�m'���o�t��(�b�!������ܑh�����^��5�6"���E-u�E�,c����+���P��3�f�����m��W+�$���M9�ݭ2.��T 5��>-V���|;=P/�l���(TG�Q3
�nl���E�6�Im�&H�!~��{�Dl���&~����(Gh�5���i�i��Lz�����%)W��q�k�C{��1mITkwjz���Ժ���̧�D�m�FmT���!g�6sMC!�DD��>�-��Ww8!�leVG�fLX�o��D%���+�C�o��p�LBJj|�ZX�AY����us���o�����צ�Ǯ`����_}E�����CGr촹.ς	���<��i
�kU1���x���1�����95y��@��7UF���N7g3 *w���C-crlX�گ�2��n������j�+Wz������qf����8����a���$$s�I;0��;ȶ�Cm	�+>��[�{���`o`�C�J��G�=?�+fd�[�T/Х��sݘ��ZʣV�f�5�*`&������ԴC6���p�A��2�hE�)l��@���3ؘ�ׄ�Y�~�_�_����U����M�Zsek���&w���:�/��N���x�bf>�Oʹ��^�+���?d�]p��=γ���)��-�ǫY��=�5��gf�Xҗ��Jzo���b�t�~=����I��]_%��!d�� �{�i.dF�%��E:w��;=I	�8�ngh���_��D��:#�k���@n�ū��;W�Z��΋)��3�Zm��[.�3^p��۾י|��~�ɣ�hQ��u��8�h��><��&�r:��{ؘ����JL��_�R�9�蟇��Os�"ȈOk#"Z�"�����	Z�H��]�N��#ve�Է���j1�-�.��6V����>(g�.��#�׀�$�Yi\j.��:	��Ϲ�[y�Q4�[���*9�{�(�Z�B3S&���H��b`B]U H��t�mL���B��Xt�T��'��UҒ7\0�5Gzb_	�dud���ך#��6i��	jQ��=�?��������R זOOG�������������l�����c�@���v�+��U���,�m:i�y���q)�#A���1��hɞ�w�Z�z���f��~u	D�m=���N'h��-ى��a����h�����=�P/Y�z�-+�T;Wv��)�g��,��]��
�#S���6h:B��zKwK�9��YGc��|�;��:&���9������!M��{́޽ő��c{${r�3ߧY$ۓ��sV[P�K��Sݖf�W=��Ô���6{V���m���O�*U��Z[r���e��%�Lzyd���r"W���.$8F��q�ٟ����K�wY�ҙ.O���x ��)��V[�/�>��wF�S�?ASV�*<�,�6���ӝ�^�9�;M�Kľvf����H������Iݹj�o��[�~�5l���u������u��mݛb���_���kFIU<�r1b�a�<`��4�����|��j�<U�VB�J8Ҽ�3�dH�U��h1�4F�zӥ���0��B I��!�h��@��6�H5Ԙ����->�*���,]����h_�u:�bu��f��}Tx�oJZ�&J'�{���ӱ��������2y���?�N���ԋV׭���#�Fj�@U���]�+a��\V���0��IɌ��$�ѳ>��@��
Nz�Nׄ��MY]�3%�ߴ�i·hA�fFFK�,�Dd���K7do1��?B�@�Ԏ��}Tx�<����`����f˟�dq!!���!7���\�X��q����3-��m��hA�Z~B�IaR�fR"ҋ2/��T?��)+�b�|����k�>��T;r���lv�B��/���`�����gk��
>��lg<e�Cr��D�V��5��E=��H;��Æ�ME,�%Ӯ�K�@�rmC,S��M��T��U���L���S�N'��㭗��&H?ܸbF�.עqz����nd�t����X�]˭.v���H ��
`1[��t-X��,p�R����K��mc�����h�(�����qZ�������_�0�@����t���rt>�LNL�f���Y����"�i�=��8怴��
�������A�Ԏ|�m�˦}���_� �X�Z���Pf����֦zi�qL=��6�<Bf�	#H��߸?(�����3VC#��~����W�S�4c�_���r��"l7c� w� �)���B��6]��B�O4bzi �4�^V��;90�~^nkb���2R�~%��b��r)��I	ڌ�os�J���M���G��d�/�T��RR�b$���
���e'�爼~��(��)&@��H��"�R�t3E.(��$�-^�&�f�����b׸��9��S�����OE�;�7��������dP��G^Wb��;>>lP]�U'	A�q����߰*�3,o7�C�ۗ��26�$�%��k�9I���?�a�2v�)}������}�������땀N���bG�}�
���`�A9���.D0)[� ���~)�X�/�&Y�s ?�~��+�X����$�)";*�#���lW��7�`�y�:i��U^I9,�S��<�ɒ�p�/^�Xb��'��ns|]jO�0&�$ ��eۖݻ��4���D:��� ����u�u���B�؏����\��^��%#Sdb��Zo#0�G"��k0>�Ƿ�,w��0���s��c����fסdpc�/"����\9�6_T	E���q��3�gU(k����"ϮV���YJZ���2sT�C�|��[�����x���xց�� A�!�y�����9��LFԚ$Kp6.�ޡ$����*y�)R�znIێ��;��ib��v�~�9^t���{�Os3��D�*�$��)#�T`���sF$.�#Z�zW�H����8	=ذ�)�_ �K�?�n���l���\s��r�.c)H��Rﲧa���^��2ig���'��f�ң����e'�;P�їd����v�_���Wv��+���6
�S��&�Q������?�4:P�ΑIEl�	����>X��վ������=��Y�4A/��63����3�*9��C���\�� D �#8f$����
��޵w��\�ztG�)�e ���f�M�P<]*���:���8���m��̊�o��O����1�K��O�q-��i��#U��S����p!���_�Ut�/����̍�"h��!������}p��}�b�Z��'���d)��@��n<3
�~̟�3�ʲ�j}��Uo:�[6�����l��6�O����vB���H!�w�5��s�΃@���.��!t��ￃ<;0��l՝*Wt�S7u|�1�:l.�́axd#�ɢ�&�c�{��?����7�6`V��㚑�����o��8V��q6�W?`��eWd���P���꛺Q�Oħ�����q�0�� T�k�8��{xMk`�@3H������C��ͷ�}���
��-"����CJX����R��X��n����?��mo�b��8��#k+ip~~����}��K�a�QE�s>!�<A��*�_�F�{S��N�9�x��ÿ��s�4��rp/ԙ	ˎ����Zj+�i�Z�����ڒbJb��\&ݜ���X:��agG�E=ݗ���z��f<��~�I���mc~�"��������ZIh��%�w�zp�_�>t��K�����A��۪��T7���ʹ@�������cF�nݥ��d�^%�I�K�l^�|��D��d�U�BZ��:�|�[w�A���Y"�q�H�5Kr�����t2���c���pQ�2_��n�턘7#ݶruu(��v�ǉ����o_P����%��D���:n�8�p_2(k*��w\�I��_E��A' �矛D�:y����+b9��[�gLFG�U�4S���!�n��M���A�SY�����KǚO?���ki`���s���Xg�@C�������8��Up)E�ӵrhp�J9A�4�����_t��6�M+{'{����o���&Ã����6;�X���5��I
�c����ik/�ȓXdY��I����8���Cz����� ~�Ҽ�Q�N6��j(�D�~ن�4��Ґ7_O�/��{��ap��\-v�=4ۚ4��Z%�}�`Jw�����\�W�s~��S�frٌ=��Zn��q��.���6���b���QRn�?�p��>�0n�����bj�q~�
S��^1���l=��D`s�����&x7�%ν.�
���4y|N~!��4�� ��M��QeoQ�p~�{Alk���	�MX 1��v��`���H>�G������yԅA��zgpu�b!��b��22Ys�.q,LH	��@��QG�0E�Pt^�ӵ�k�=DN�,��T���恑���T�z7�~�}F"EP!.�O2��TƕHW7k����1-�c���~W�A��N]�;w<A3�	$�)�
 H����#�1��������bR���~33�4C7)��}[��_.. ,�D�^@� n������'�<�u�������߮^�$7U�Ys���ϐ��3�[���=�i6=������l�F��)BPWZ���~)�����?l��%�4�|�V�I o�9ߢV���b�
��i��3J5�^���KZy����HV@����-n��3��q�p�±����7g�CW�ޔ5J�Dg?�o�7ۤ�_����.(�����Oګ��K�a@F�+b�tI��L�z�G'��i#4�xkύ�E�R�ã�N5y]VG��J�N��S�_ ���a���7a�*΋3C��,J�ښR,�s�y�]@0��o��_�G��Tp�:���3����׾�&���[�wr�T�: ���-��S��_c�1�ҷ�o�<h����+�9�Q�r�PP�B�9���S&�ﻚ�&cr�-��O@K遬��j9O�=[?�j��	���q���3�eTgk�Ii�kl7��hg�q)~�y4�����i7�HS$4&_�C}�����F�w�*Vș9�e��{Z��V�������^g�%��i�&�Ǣ\��s�E����������%'�gsJ�5�/��z������5&aIQ1���>�5UP_݈Wj���o������r�	��t~������Ҽ���c^��b.�GU)�$�͛Sa�r7(�K�n[���'s�o�_�w�F�L�`������h���V%�!���y��?�I"�\,���{T��Rz9�V��o�-��q��t=��&��jm��k���&�H�<۷Mt�lA�q`����y���p����\�z���3����\������l���w�Ŕ{�RtmBV�ƾ���k�ə���:P�2�A�~J:j}_��d�;��������>�'�A �h�bss�q	�~�2k���2���]��3W[�n��<��z/���0�d1a���|h�]ck�o���y��-�K��`������&�J0�
�5!T#�)��9y��N��ɭC�dHs𻥩'�GL�Jc�����ip��cB�\(��#q#�mi��J!�qԻ�hW������U�0C��o�N�����y�o��O4�},ú>�d�Ȃ���z�yQ��L�<9��oK]>j9o"�rm����EJ�O�ޝ11����oe�����`u�OaBY��us���văl^�1a,
�<h��k���y|yDA~���%�ON��n:�ݵ+��mܨ��|fȃ�K�s���f�֘N�MY��%]$!W�?,BÜ���z+�feMm=��)z���?W�%<X߭�����%���gCC��;�wT�ؾl.0��P��k+<�l�PY����P� ��Z�G�7I�<�[�:�`�t���5c�}�4c?U������2���sD���㕪�[�QC}ݨ�3�G^R{��ͫ���r�֗�X?2���[�#8��M�뉞ku�k�wܑT�Ft�]��vmJ>~�J
v��^�<Y�IԄև�̪�H���ɟ��ƫt<6�����5ײe����3A0PW�F�Ҝ��2�^Dq)Tt����eI�X�(#g@<�m���QR11m[�N>�7�BJ��n�"E��T<m��c���S�Qb9`����O��LM�I��I�A���0�Q�����i�/��k{��2j������6X�Et)�kW|a�Ý�������{�ڔ2B����#���N�8Bv�n (�i�_�����Q2ޟgq��HB����պ��'dD��U���'c䃙�a�=��򺅘sª�2ƌ�M��h��Q�s�Q���-��:#���sE�����q��O%.�Y֧~l��1�0�#=���WD�{�v�::�m�>:*�sIm�&%�!��-�%��YN�!�t�����H�mWTeqr4[�K�Rq���WL�=x�VV�6	t4����n
��[l��Fv8z�Q�?���5�M_�=���%�Wr��҆k����#�l�(�Y	.�ӷ��1`!���b�H/��e�m��/%��֧>���L��E?�W�,ζ��7�BS]�4L8�Xtٚ�,,�T6�q>`�w�n�HB�����ș�/]��[��w=�-�~N��ri�#o��q�]�e���E>��(�<���^��c|��k��w!ۿ��;T��s:i���5i�l�/���ɺ��u,�xu-����<M�2�z�ɏ�%��Y��7�P%�>�ӑ��B[U��9�����`V�3s�$s�o���w#�$䣐�,�׻6��Y'\!� ϊO�-���y>��w�U���G�D��[]�_RK
�)�ӥf�f�FP�,�?���6��x,�܈ <��&4�E�k7��jx�.k�@�&��#����ՙ<&M-��w�cK�>�3Y����`w�6C>}�a����ugv�.`����P��w}�)�˃O�Bv�tͬ��������_�ɺ'����A�:��o�y��NeE���T݀�S5X��ƻ����iƾfu~�@�����<u������2IKK��_���{mB{�6��x���~��k�
�� ��5�.<r;=��&��:Y��9��I�x����CnR+E�m�61���������%��\�v�������U1s� P���8U�[��q������~/�������Njdo�g��8<��SB�r���{��@[���� ����?���j�X�i��z�kt�_������
���teC�#[�7S���1��O�|�S&x1jm�c�yZ������Q��B�3 G�OA;�����X�$�hJ����T� �z�V&��9���Q8&��1�:P�p���Z�<v��t>�7��]ko�'�RjBi�u<�E����l���
٦B�Ts
���^=�=jM��v�����;zbd+�lJ]����s~�I��~.V�k��+�Ԛ�l7�\3����.c�<�9���0x���qŜ�����x:/�r+���%y�.���ￕ&�R�ؒrr��,,�QѨںڒZ|���U���c<�ؚ���З8�^�e�[��p�Ѷ���5fE�e�����卜N!3�t!vQ�`pW �֏����S�,��Ʌ%������h�KK�_h�R1�ejVo�<O���t߹\/yX�M���loE[�s����R:�n2�5����
�Ey*�.3=��y��Yjj��diT�[��"pQ��3���6�z��T^�RG�E&��d��N�V���j�è�Jo���bs� 1�7~��7�ـ�69N2��n}�ʠP�H$/�ī���ɽ�h9<P��n|���ooK�V���	Yuݹ�V�o��LE� e0n�7�18�k�*Gp�t��PA>?\y���m�9�Fl㑗�C)���q��"2t��Xb���i�=|ﶶə�P��#I�I*81������N�����}��F29�t�W �bb6�vr�>o��> /�j����!݇���]�].�HBw?{�.�^����0�?�9������Zym\�ڳ�0A��+�hȠk�����j���M<�[l�i� �G�<ې� ��_	���xT5��H�X������0؅)��}I%�yGKK��T���/�R��,)f��1�e�r|f���L�IC.~I�$k��O�����rG�����$D-���B�h(�Dml������R�=X�eqab=���[z���n���}��pX�+~��x��������j'/D�q��R��7f��M��)���G��f�g�s�ޅ���=۷}��G�	}_~��`��BZ����t��,?v�ɷ1`BR�.Nsg�˘r� )����~����3}��_տ�vj�E��Vw�и�^�z��FI��:�0zO�,�z"u���hn$�ĿQ ��cQ�+a[[������}�[J����H������р�c���{�ِy�3�����L����`٢���I��)�ZѶ-z��o����^����ң��·
��Dc�e�TD��j�Q-��H-�؏��j����Qo@u���'W��D�k��Pj�R԰�������a����(�C��Ad��w���j��xQH�U��RDj��*@�\J�tn�}2fD���WXI���+�>^K8��9Ҙ�5̫bb�@dK�%���A��I{��!�h��8��ډd|�dۉ�%����$H�nԵ6Y���m:k�:r������ى`��s~�Dy�W*2�Y��U?"C�B����+m!Q��nnn���b�w�e��Eߛ��[���ܽ���	D|9=$6���~�������+OG{3a6�9 �ؿ�s���<�:���1yvs۠�䁈a1�4�����a0Tb+�D��	·� ģ���}U�#����éA���r؄�O´Ԥ\]y^:�v��r�py_k3IK&��E���:V"߁f:�%���z�LD�Uj&M���6�>���f�k��nsU�Ƭ��Y�� y�@�#������%֣*��6�vB�����N�֚�+��������9��� �F�-P�� �@O�0��ӓ��Cqa��H�A�ȄM�]�E�RO��[>��k�R���f�Z5<��p��B4T��IH<`Pe��{G �vDX�jwEA~��{�ܑ�J_u�;���0X2�>��X��D(^A^(�ݩ��闫FF���Y�M��x��?�~��	łY�kD"���y钥Jl��\���)B
LG2��)��'0^��j�x�G8P��Ҧ}28v����1�{A����IFJ�T���@BBZ۹�^���4���� ���p"ŵ� -��T����!����~�>|47UI,�m	�C����|���$� G�m���>��;��XF��S*�������&�У��� ������]���!�?����EoVC<w�<Z��5���ns/��г�����*+��{TM���K�+�z&�����'h�l���:����&���_u�1;���2����Q�}2�@C5@瞴���k쨨���),�C��:�~qqaz2��;��� ԙ546Z�}%��m����mhj2�.Q�m��5���@��c�0R�+$�W�� 2ۏ��oн ���`�\��|9�BOW�t�m�ԭ�EG|�jʔ
�X�M+�� ����f���^�ڬ�e��W���L�+��XR��zH�h�=�'5c�{9�����A��[���E{
9�"8�a�/���.�̨�*�؏f���H��,,���=:)�:��KR�̩+��]7�SVs�5ɬ�����W���;�Oe�#M���W�-��k���BLPo9��{Y'Xq��8K�;�-��pZ[O��8�^�����-�|����	ψ���H�~�ֿ�ϙ_���!�r�{�6 eˁ�0`�I�к!������թl�h��������3�5���+�����s�������Q7Sm/U}y��t�Q��UPh��[b}�u�����w[e✝wTj�"��Gߢ--K�9^K�V{O{�C�>/C%���v&A��.�R�$ta�a.��Xr���
j�Z"����(�j�������k���i��֥*Z[[[/G��X��CD	�~u(��s},��*a͚��G$L�7��Ԃ[�l>;g(`��bw����֔����y,r`����1���\����y���<�ix��M����+��nŮ��d����Y��+����ى!�h>�Ǽ.���@�]��g|NN�K��"�UTa�6�AhE��
#�hDe #K��}G�t5d�}���R��[�Q݁����G�1c(a$l�9�ts1/�����l�[��||w^�'����p���p((�]��,x, �99�hk"}�U'@����t��&(�E���ϖ��88��uk2.Կ��:,baa��:���� R]����"�����Q���n:� �t"ZՉt�'C2ЇP��ֶ�8�G!��R��lmp[O��� ������o݃i�A��:{�6��cҤ������P���nӐ|۽��Rot; �*�@I��Ҥ��!ߓ�j4�o5vKQYd�M��,W��ӓD]E�7���}�-�����#b.��g�4�).�M��:�FB�D���±�Q������6��ѳ`q�QPJ'�~~J�{�=��3�b"�=nLs���<8.i)�DO�9� ݎ
er�]>��[�,�B��#��o�[.w��;�����$�ߟ�f��E5�a�G�-�m���)��~����}?�|IWz$j={�_VZ��Z9����N��5o>���@��]&��6q�%$�;��vt�uIc���d��0��cg�x�#�|����mh���z�bd�Uo�F&����,�LČ�P�`k5���SmG���ҟ՝Phjz:��d�/���0����t$�����KY{049��_aޒ�'�'�xOw4��Ki������`����r iU�&�+G1W����U����� �+�e�܋���cQ	��Hb���.wG8�?�­5D.[�b�B���s��Ė�Ի����W�W��@퀖zk��N٠�o_(��g�(��g�{�3��A�6,��8V�8DA�\
��G���]<�]����	�p�\A�f��~������^����;��@��Zw@,Byhd����nt]	�IrugN��tS`C�x��gY��2,cbz�u�����ܳ�yKI�:x8�vg��V���'79�B(6�XI^upu�Ĩ Гk���>X`Bp��C�2�Á���K��5�����D]2�RM��u�J��<�1�f�aw�� �S���kg�'`_�nu&��e)�/�U���GH�iao�!-�&��_��)���h�q#��BgCl�	��
��@r<zy���Ef{L����ME�Ҹq�K�,�䞣w��]F^E�(�U�b�𤋮���Í`��`�����|��������&Я��0c��2��3����}*n���K���[��x��WРұ_4O@#��ӊz��S^�5 P�j��CD3=�;Cz���*�xߪVM4P���np�Bq��O�u��)/�)OT�f|�@�R���-Jv=�v#d�pW�� � %?/�VA�u�.����&�$�`��#D3�P��t��㊄��B�1�����́�K����y����/AaYș8;�<��[C���{|�uύ���x����l��r./��H.2�$M^���}�Ŝj��ٶ}�IYv�E:k7ϳ?⒱�)�id�~�������/���lm��`
z������q�} ��8���u�Y�o,}"4AU��*��Yn��,6��^ɩY"�^D�3�Q7W߄.���9.J��Fs6~��:j����UV���V���[+��ot��m:�W��M��<�E띉�b/�I�S;#�J�� ��\�B�<'�A�ir��Na�����煉l�K���ިפ`Ѓ�U%BvE���`,�8n�W��#
߻�RO��)��H���y���ђ]Z�t����n-��w��)2��W?��A��'����^�Df�����vh���P��K��λf`wЉ0ܵ�
�=Rts��2a�r�g6�ϓ5AB���6��N�	b��B����r�n����/7NMvH�@&}�lL_���(�
�v�-��2���L���]5̿bDV�]�_Q��с^Ŗ%X�	91J,I����Ә��_Ϳ,�X��*�![P鉒�t<���gy���|��Y�s���(a2jh���9( ������M]4A��B��s GuǗe$�~��ٟ����#�.��c�$Q�O��"��:e��ۍ��;�M'���+�+�wگ�yZ���&�|��X8�_䉼~��ް�v��xTn�3�[9hq6�̇��r���� '��X��I�L���W�!�SDJ?ck�	mS��\�r�[�z���(���eu����AFLr���k���[X=�q�0ø�c��H^�v3=^��<hĘ"*A����Y��_4��%y�)���L�*�q�m��}�n�+\�F�����Յ�|Y�k�(��n"�Q�Au'E�)�$ "w[W%�8u�����Xf������LIG�WM�/�#'Q�ۊ��)D�� ��\|�7�T�߬����r���L��>�,y�m�Bs���Z�L>k~l���oL݆�6�@�9�~���Bd�gu�q�l�c:���3�j�m�c�ms�QLKo�����'��&鹫��O��"�u��W7�ޒ
�3!��U����`P����$(�ԉx�򡨵
�mvN��:��͸;��~�~��@��W`���t��W
��.���E� �
&��G�������:���vG��u�U��P!Q�ޤ1M)!(��@���Ӱi�>Z����D|�_�Uݵ1�2���і5�&����]�}�+>�.ح9���:��N+�Ԍ����x����p���ʐE�7������P|�8;�\�=���0����	���Y�������3P��VÞN�k�N��K���F�W!zЈ��:8`U>^����|��9913�e���~t��%���R��J�|�] �u�P��ر{�������� �����C�in}mG��������y���/R�2�_��>},+���Q_�#������N���j���h�[LbI;����݃2�u�4Jo�nsʜϭ���ytk��q��g����7p�xU�,k�%'����R�%(^nJKy�	4�1}Y|HZ)WM����n����@.]Q�"2��Դ����=:�LI
�����^!z�~R�̟"V|���U�.grwv��8,X����?����ִN���[���$ʒ�H�yR׽�`53�����5�p�ӓ|7�s��z�m�����i��p�`�g�U�|Q��0�8�@�c'�F�o5����pWӑ?'��]hO�Tg�����1Ϯ?���0��޴~7�h|q[s����m'�p9�l|������k6fV�3����h�A�T�&)���`�	��f�ۣ��$�IcL����:0ȷ[e�Ź����0A� l٘;W���n� F���]Ȋ+�����<��v��Xw�R�J��SB��	R�s@K�]��'�~�T�H���]�Ϣv�d-C�.��j����j��k���}�_��Ү`G� dac!:��XTB�?�ţ�Uh3��9N�5D��=&��/������-}<�5�Zc<��9�*)a�v�_gQ�쁩�ǁ�#���icJ����$�"o~�����~=��̡����!<`cv`�z��?��"�X_U61^:��w/5�:��y��֊���tл�z��朊#oo�ɖ��86�\��0���V��C�wF޵С�D������yk52���:�����*��1	bB�S"h����zI�P[iO�����E�D���/(a���w��Ƭ�g��tl�Ӎ����Y���ϑzH:W��6T\}	"�Y_PR�����)�g{����AtA���U[W׼?ՖHScW������xU�.�	�<o���
I�ֈ��**��t�~-��8ώ�
���� ��Wf�c��n�4=��"���*XF�u����[�$����~��\j��!j���TLd���(��R2���΂�~��ɉX	�t1[_'�^(�P�M�Dރn�)܁�{�Cz���`�$Cm-��TW\�8�z�16��!�Ђ��Qv앸��"�W��,nn˝�A	��OClՌ6���XȺ�=4�q��x�i��ZΈ���:-���(H|}�*K��l�a؄��1�((�-e�~�7���%�	�:����@�Tc���8h�7���E�lXz�
���r�Y�8f��+1��n�O�$2D��~� �|�/��p��K�CJ21_�1����rs��^q
��Pj;����j`�_��닉�E�G�i%
hd�uƐ�	��H��蹜����-���Ⱦ���Ͻ�jW/�}��oNܙ3�N�7�ĥ�$o�,o>\>E2���[�Aq�0$3��Ǒ��1WZt�I̋�3K��|�>6]>��=���Cw��&^���ZT��?�H��Y"����S����]�7Jns�+��C�-�6A�'��FF��%�f�ݏÐ��P����W;T%���B4�:���Eo�'�_�?�.还��~����r�1(���ɻ?='�����dm�;���U�lY[�����m�?	1��G6~��*z��o�[�}���pq376��1Ŗ�ª����"��!M
X�E~D���Z�e)�y//j��/ו�i�U��ݲ�jH�Ռn����P8��M��ʪ����'�כ1��*1���A��=�4ڦ2���j�F�}02�7_g���u�����ii>(�rO���0�)ҽ����9�&k�fub�ڠ�8H���ᜅ�,���Аt���5����A�JNx4�J����)��r���Y1]���va���Fp��A�<	))ࠪy�A�6JG����w� ����rl�MlUVxx|�)]_p�?�U���!}���W�]~R���@�7a>�T;_zQ�Y�2��.�?�_��������Ø��z�&q/p��M�Z�h���tTP&0`�q�n�9�.|���� �:P�$�N9n:>���`v��0�W��B��Q�[Z�y�
k��y!Wf}u���8�馉s�
� } 1��ݽ=)y�c���"����EL�Z|�,XP.7~�Gy�q�gu9s���u���7#����H�-^�O�������s8�o��$��!f5��qyh,��a���W0�+��M��R���I���K���T��ddrKKb6���CE"i-�]B�0�4�B�/4�{,�E�P(��O�X�Y���Gya�	�U�nK�c��ۇ���,���I��ek��Զ���+�E�'�$$�G�����|��8���7�W���9�,�hi�䷥qh�HnӪWgs�>6,�ik��[d�,�cHNC�rG��z4�DTa���OX�S_(
j+��"=<]UD3K6��{�ַ�?ؘ���Uڃ<$b�2|�-"�6;��,�KW}#��C$�Ϋ[�0F���q��P���-'�{�)�NA�yE&ވ�V�b
��)���6��R�6t�<Utii�����Z�t�!�O��{��ق�����&c"����Z.t_8������aV7�GS�(��,fTo@<�l�Qz���K�����:�f�S�ӛ��jE����հ��1�㎈
�|� {�m2��,Q��4�H�0���xi��+�f��1cϣ,�GU�uڼ��� -�F�;<�I���7���v��Q�/�Tک堫٦î��#�q� CA,1�~�B����%�a�>����؍ ����'yT�[A��"p=���ewW�r+�I�6TR�
)Z'+���b�����K��q�8�
K,8�t�V�A>�wz:J��	�82�r��q��m_#hҙOA�����;��k�d��F�[8���
��޶����>)x� 3�]��ǿ���>�>�S	v������LN�П9�aV�	����:�̃`�%FW����4AGG����aO6��r�	$aџ��}۷h��NR:˵Qk+T������ފ�u����c�T�Z��Qt�0ij�l�w2vv�e�WėY¹�)��H������i� �3s����Hc��f9>�#
���A��/�L2�C���q,L�);�c̉����@GC;�E�����j,�����M7eU������6��}�m>�z�r ٛ��[�E1�a&<�?��:*�����S:��S�.I��隡�SD�AA��ia�!��!���{���5���ଳ�����s,���·�ArA�7A�?ҏ��k��F�X��T����'d�Þ��n����]]</SLL��Ŭ�$��o�&����i���[Wv�"�Q�d=K�
 ���/݂�1�ۼ:|[ǥ��W�v2u����u9Y��u���w=�vࡪ�W?^EU���'Yk-��\]��sw�Z�x�|�@�����;{Z':R��~?$?�JKKN����P�@u�޼+���k7b���#�h���OMV��g���}�viݧQ���@1Gl�0���-��ڮ���L�&;	_��p�nl?Y��-�]��/Fŗ�������s��OKio�U�;��Z}8�k�gn�ך~���DZ�h���j��*EHb

�u4I�c�&��׳�lmK]��gA|�+��BGG�ւ=r�9�GE������3;4E�f�ŕ��ۿ����1�ϑ��$����������_
!��&���Fh�Pq�R)�l0���Z�u�⽞pu��x 	UaN�ñ�WN�$rZN�:V��y �p�!�ig!�0���G��*���Δ�јe�ϞKp�͇/I�d�c;��	bEU��R{�C�kB5�Zx�Z:��ӌ��v�������-��.�V�B����"�u��9>a�zZl��{:�-��F��Ġ==���.������]�YI�?�����Djk�>'�@/��ʂ	v��/�����X��U
���;��I�0Zt6�}��w-�dq0���m���/�ϛ}ha�4sE�Eg���V_.$�4٦��_��*1[�=�o�Q��>���c��P.W����yj�2�NVv���b���Y�W�/"E<���L��&4p�w���|�L�Th=��!��C<�@ ?��4I)�i�r@�Ԋm�}��{��� ��f1 �d�$D�~����H�?&���,�$����Í�d4ùJ� #��-��E�?JNK�Wd�s�G!��ݫY�[ſ�Ԛ�����fP�LS�D|�}M/r*�Z�uw���v��X�ť�njW�Ly�Z̨����¸���紲4�ӑ�"�vg��|��e���L���Svb�߆W���WP��oT+��0rj�*kj��!����[�����A0�i��N�Z����;�^[��Gi�N��&雗�~�T�ߧ$�>\cz~l�lזy5_��w���	w��9��.S�x�$4�~E�Qa
�r>��h�4��܅�K�*^b��d�?8��Tֶ����d>���8�&��3�>��2W��vvj�Xp�!>ٌ-�oO���'���a%���10��AW��$ؓ[ �,����%��J7[t���c�YAi��f
+(�*��xr���6&C'�)nw�}^�������k�$��_2$�=�%U�������1�;�1h��˪G�O!fy�-Tn?�c�&�&��c����6��r��)_�hSK�s����Aw�䃣_�xS���x�˵B��k6�3wyRHn�^��p����^�����u�'��5�K3����+��;k:S�;?nV�X�fB�����S��90�Ԓw�@17�t���^�fg�{D�n40'����WVjv�BFh(:#���$�A�:��ظpwC'2cu��̚沉����&q>�`�JAj¤��F
������ �9�	n�$v��g"m��=+ޏm�+s�������+��OE�W�j��0g�WQz,*��b�ϕN��
�ʰI�
w���G����gffĭ�h��^�9%#��)���J�=�f�N��6C��d���?�����E�;̐+�� ���4�8	��3�C8Ҳ;����F|���3[(ޟ\������g������c��^���.����\�=��[�rov���(�����Au)��6�d�Z��N)� 7MCl��� S0%�Ve,���:�Y��sa��3��L���{&��ߌ��{v 1q��ʼ�fܴ�]A��4>ԉB��r������	�	��Α��>�k�6��f�&���^��:���V�_��Yd���h�v��N�~�6�da+�j��.o�����E��+v���k��Si�8�r�К�P#�������r���+�Y�g_���[���Q;ntJ�g�)?�gǵ�Y�.v��c}�C|��ɕ /Z$�Ci��lz@A!c�����{՞ns�r%T1��״��pW36��<�g\IҼ3u���t̃�t�����L]ڰQ2�ݘe!v�\s`k)���(9l�Z6Y��(?ں����iZ�����Z�7�Gd�}�ж���JM{�y�'�D���"��=�\��f�`[k����{��W�Y�<U�D�~�������z6,����n3��� A�[؅<7�+�ܕ��=[�
��<�ʥ���y�*���i�Eȗ�zng���g�#l�pz�2�1:Q�$aX'Κp�k���=±�΢ҍj���U�P�� +?,w�!�ɋZ_�����N�����	�.���n�W����4�����2���>��\����=Wx��FQѹ��hv� �<�6+I�a'U���,��g�sav"���{F\��b?�*��{����[�GY�e��pw�����1���n��N�տj�-jƂ�:���-1�1E�G	�ÁQ���e����ʆ�w/�-��0�q���V���:wa��g�|����y����-̰r���t���`؅FXy�3�����sЧ��[�;��X��Hk\�c��>�<=ۭ-uA�1�I�J�x5�a!U���՛{^�Y�e�3I=�w*��.��i�?λ�Af/QY�7�%3~���yv5I�[W\G�$s����4�~�RWUH��0�
WCZ����G�������̆[Ƨ���	�[i�-n�GxD�n�*��<u�H�5�\�;�\	�{�z�O-6Em��j8��i��ꍍ��7Ű���͐�����E".�Ń�:TdCqdy�����9�2,����'_uǿ�TT�H.����_�+����}��Ӭ��_B�յ��4"Ʋ���"gB],1���x�'����)� ��u���)͹�Dϓ�5Ӭ\]�KO����%�YM[�3�	��)G��:J���p��L:��%�c���Q5"�9w<�R7A����xn٢����"��+Ո���5f���@�8B(b�2���p����6�o4���\���@̪��/���<����f���w&����a+}�h�ڔ�m_r�I��t�%��3hG�d�Z��u�p�˩�2��#��ۻK K�>�qK;�D��&�i#$�E����V߭�'��*��*�"-���h��t�A$�pC>eU����p��Ap*�{)����2W���*q���3ޟF7[?�O	�C]\j��t=��6����ͫ�����X^k*Ə���,��\'c���B��M|��ZJ���`as���'\�nwvb�F��/<e��A:��cU@�2��=/�g�x��~2��8�ֱ:a}J8��g�$��)�����m��,V
��2}�'���b��@=��om}Z��έF��F156�[-'�������}2h\��?١�O�00���g7���!�5����u��b��)�+�$C��c������ȓ�� �ZD�
�#�g����Fr/��u���(T�:����s�p�[����ëa,����E�q�7�$0j�p��H����
�Ȼ��OZ/�v�*W�^��5�[�B���	�6���"z��cR�1��XB������j��l�<�� k�/l|�t#��W�͎�,nV�y*�
4�Xlۢ�$��U�m��}MC����_\Ot��������>��g�`���b����_ʋ�\�ܸ�ǯ?��Hx�Ny?dڞ��Wu�|�Pc%��F��;f��.E��ty'�Ɔ����|D�M:�㔗�_�e����$�I��+���,���̾s�p���e�k�$:|LT�C�K�)��������o��.�| �flՄ�29o7��Il�����s�Ћ�d���zM��R���?k9�'ö͘�$����M�5i����[�����'�?�@}��m�w���K�lbkŹ�w�l.�'�A�W�?�S���>�?�2���0^<���%E:O�뭁'�Q\%�%��j���x"�R{�a��w)��l�.�3=ny_��H��	\�Sz�����7��Ч˳��\���,��Tm��f,���V��M2g�p2[�'�������
�N���Ob�/��C�/����k�3����>xŖ�3���(����e�����6�3{4J�/��h�iDy_��ʈ���W5��9�X���D��7��2_��h��@;�hh�9�*	`E��@�X�|�H֣��+M���1n0��͹�H�|�E(1���v�����n~��D�m��Ʊ�4�;�y�>Kt1N�n����=+��Ý�e%Ohбw�vk�Ѐ7�b�b�(�򂶵RYScH�Ϯ��	Q�p��#�zV|ZVܼ�;Z�`�+*�F�ɩ|�%Xd��;L�����ӵ(�! �vM}X���\��X��yJ�����u8���6-_��x��s���4�D����[��1'����hc��%�ធ���&�3d�sx�1�W̧�) Q~F�V���m�7����ϕ�_�d���_���z3N����v����q�s�-�V���d���g�+jڋ"ĕ���=h%� ��B�A����G��������HG��v�5yq�-7���B��r���9�I����)j�l&����	ξ�P/���C΁�sXP��ŖI��E��9��2�%'��`v7H_V�{ǅ�w�L�*�Ɣ�>�t�<K��g�uq��*nr8"}�~�{+\es12��T�I�8�����8���qI�Ut��#+�5�y�wv��k��0�O.�n���V��l�//.e�r�������r�$�Ɨ{�!��h��.{�G���r��?�]ޣ��9[�Ns�[�_����);�:,��j�4��T��~twy��ΐ?�a�r�t|t*��{<ud ���t���]�n����E Ua�_1	�C)ف�b��]�Y���n��XMw{��å��\��J�~����$S��eEf���9�S�ɗ�M���/�>�I^)#gI���=)p�]DRyV���sW�ĩ�q�IasZ���u.�Z��a��X���Ј���c|�b�O��K7*性��e�Ҿ,k�0䚥�|A�Ҙˍ�}�KU�t��m���C�KЭ)I�'�5W�}�s���9 ���=���[!`�7fA	����*�`l2��T-~<F�_Fh0���%#)�Ά�Å16v��w�������D�Ify�C~�1�JxR��I$T��	���<3zv�G��������ox,��{pPna����5p�υ���ur���AXK^ل4V8@��79�B�X�&^���_PV�ۥ�9;��&�Kc�'������S��Y��\����jc�*I0+3V��g�j��K�g��]8!B�E�	p�7�m��<Ί~zlɾ�5-�d	����O�YvM�>�f����靆�Ew��[ޭvܲ�-WbouZޕ�q���%� nWҬѽWW�������,I��w�Kw 9��=��[��2'�xbdϑ�������* ��� ����������U�c��IeKO�|BN <�4���q����L\��T����2�~����^8�q�.RV[�<���]`!E=� �N�_�$�[���,������	<���ht/`'���e������R[�1�-��o�"*�N�k��+���ٓp�D��M��ɕ�#�g����vY�VW�D�����Y���M�B�$��W����>w�a�(���T/@`���B�84gزeTΑ�K-��.ǃ=
��c�pT���vt\1���5�g]�������G\�� �}7(7���̅	�n���"�9��/��ik�/&!`Ӻ,���,v�����8ƍ�q�>C�'��Z��P�����J	�zG�?ˁ"�Ν�#��9-�-��R+�a.G�}3��2u8��9�b�_	[�p�8�H��-�[�C^���nX3+��9Q�O�o1G=w�J��[�F i����~���PB����8��F5�V~�:�b�t��Y���e��*+������Љ�Y���=^����`V�O	��+��X���
+�]$l�d�������� �� ���Ȝw;�pI�u�7U7�Hw��{�?�Q�ʬ[���/ex�����q�� W�vؽ��&<z�o���ۚv�[=�K]�]�@���Eӽ�_^�<��>T<w\b�@6HÍ/�I�V�F���KGW��6~�����hi�*	\��u���uM���Ž�;��4_�Km�XMz|�)[�[nN{���O���i+�/z^"a��~d��L���#ٺ�iC�}o�<�-�W�N��;8�}U�ÅS�����7�3(1�z#� -�����p$W��.�����H�AK��Mn�`��bO�4�1��ٿ�5������d������p�4s���Ɖ5��c��X{�Fi�cc{�:�B�{�fc���[ �p�,ꅘ�G��L�W��	~k7��|ςڿ�5~��~i��D��������Q��2q���mA�Y�Wl���ӳ]}���(�)���z���_W�p�IbJ���U���U�}q�U0/�n �K��O�/�e������zl6�n`	N �iE�03�@r.�Pd�+�b��í������e�5}�ajby��z��!�t|u�	0�+\�ѧ�~u��eV��i�3��ox��(=��V�o��Vצv�f�㯱Ʊ1���6qS���k�h�� �+\nmq�r3���/�d`������[���ڱ���B$���~��k�Bx��
Z��źZu�W3�r���σ�m?��Pj�=[;۝nv]{>[e����f;I��V��4b2g�U�`M���&�ľ[Dk�����d$�M-������A �\�����ѷe��证j$���^��gU�&� !�&���Dk�@��}D��ٞ�UبF��!�Ƨ����m��	�sL[��H��I��W��Y�����*EA�X*5�a��{��u�;aϋ3�|ˮ�&|��r��HD
�k�fp1M����4�,W泛��&)�Z��;nEn�,�­����	̺�I�6&S��	�gA�D+5������rL�mv��5�|Y�_{\��A�s���^�gG��h��}P�]�W8���Ջ�5�*��-��'���.��Z���s �S����Stt7�;A$#��&�u�G���[��}HT���(�!L�e/Z����H�_��{���%ԇ5N���W�IyI��)Z���O��J�b��>��������R�K������\Hn���z���G�}E�ihf	��	ש��="�p�Bu��B��]�pX]�y8v�/�A�@����X'�M^:Z�r��*f�T5�@f4��!�y����d(�LĢ`��a�k��b�+��%�+Q\DfT�e>.{?͂�
0ک��J���x����8�ؚ��3*cć[c��?�A*)�����a�������6���y�A����zE<i��U70!��I���!4�Hw��4��ݣ�;���;AGN�ֶ��M�ogg���X%955����g�(�x���0��q��冱8X�z��f��{r�>_��Ķ�1��y�m�`a�9��lH�8D[ϓ/mh{>�$�����ً���Lq^��ǒ�t��:��.�3�d�Ę?�K�YU����ԄҮ��'K�'�����-�5�D�}
�t�pC�'M�0@�"ڟ�U@\$~EĬυ��&W�b�����Zwor�_����a.{,�z���zmXJ��,��x�˂��cr{,�()��I����}��'���[
r�OCK?Re�~���w�N��-s�X�&�8z�h�~Gơt}x?�v�wYg=�z�u�"2���%;}D��l���~2[Re�`߷�RjWjk�8�FiP�+N��5i8P���]]t<%��z�&�3�P�]�4����׋=H�֘�hW�E�c�p�/��ċ��˼��%�+;��Rlۢ��CD6�T4�2XE��o����t'��bg�h�Xl����<��J:���o�S�CI�όJ�+=V�.���Bw�b�I,O�gr���,끫ID`۟��@)�걟͹��1�[��k�u�ہq��|u��|���A�A��W�L��T<��ٟY$�B�7�ᔔwDVzuYxqx�A���dalln ���d	�'����^�-j���޺ݤL��{Pb@n\��6�Q��+e*TI�Ӓ�H/�_)����Z��p�O�����?����܈�V���b7ĵtcW�Y��6�9�Oh�2=h�u�F�a,���I�K�cZ�c5����s�I����XD�5�bHٟK���	Q�b��PA�%lXY�tg��c�S~}� ES ���#Wd	S�if�ķ����gY��I��\�
}2S�R,������P"���F�(3����m=���"���ʋ����Vg�~�{�����j��ô��?����h�"%�������Ę#TqK3�K�C��B���q�so����p����v��,��Ĭ����?+hBK����>�Y(=V��MB0��g[��r�Z�P���8�L{��|�+�'��;�98���ߣ]�3 :,��7����2��*�ڍT�	F$.J��mJ5���gJ��zpaU�zs՜��\� w��M�֥���Y���kL%]Ms�?{/t�7�Z4�K%)/��,!��|B��~�y��p�)�F+%�6z�r$��y�X�ȫ�osd��"�l���7f�V+N<&����q�q>!������*��8���1-`Kx��y�&�{�)|�g�J��-Ye�[Q�L��;K��.=�����G��$�3������
�hV��n��-������+ss��-m�o�a4����v&F<ݘ��vۍ�ia{�U)��g�	,�>D��f�
e��gPdVSp6��_���K�� �����Jf���7��� ��6N:�Pe{j�
�/�B�>��p���~�KZw4''��R%����\)�W4'~���Z�.�}���E@�_����a�=��A�k�>c[�4-n��S�؋X���{�x���a��4��"�7g8
�L��ؐ M��B[��VB��#�^��b�5�s7\�U�c��B5gDh�\2l�V��<�U�p��7��� _����*����-�m�Fs31R��5?�:`_��.Г6!#�@������u��P��xNω��$�ʸ(�E
��г���eɓ!C�"q��z�V��q���A�F�����	����?��ݒZrx3fV�s� ����5R y�@�������x,�&����Q����	5���#�~�9Ot��2��_��ܘ&��_�YG���"}�'�k������_� ���19oOv��YX4/�98
�B��g���b5fϾ���:~��9r �qB����'1�]H��b�����XLL.�9.Ķ��g:z�����L��R�}������7��4~�h�Qi���[:+�#;l
�|��q�������2}���W�c*�~Fd��5X����N�#�B,��W���~��/�����P�.��<׊�a��;XeM��6��� ���XlW0 Ӫ6��U :5����gV#h4G�!R���lc$`aʾ ���ί�u?���K%Y'$���>S �	נ䳺`ᣞڎ�`-�w;�A��v ����F@H��f?='��׆�^�sꏕF ��p�e��N��]����lWИ6Yʤ��
�@<*��ῐ���޵O:�~WR!i�1Uv��WG������ŉ�z$�n����Bj����o����!����ڔ?\�ߴ�] c�2��O�P_䌏{����ϟ]��0���W�7�����I���څ*����!�!c]���7zhl�j���	��R�A*��~m���^*�a�+��>�ja(���X��NX>�N�xb��aA�`t�.bsz�:�"����^{��;vZM_1�Ç�$�vL�� )!�yc5}��W:��c�JM�k�����VV���27�t��,[I l�sr���q3�Ek�f\���Y�?�@"�2�T$�Hbig��=���.�L9�}@-LLe�DZ��^�#��O������Ո�w��v��2� �~�:B�-3�^���!�ԕ-���`3��C�N��"tAg�A�EVY�B��ҝy2~���\�K��㱗,�0{�}���iʻ���;���2b1���G�ҿ�ʹ�8�?H�r�GM��g���	�lP�  ��/�/z��2e�^��3�$gj�K�8-�N��2.����ђ�! �(��y��&ǞN�{��7�ק>���ݍњ��[�æ]|�_�tA�����A#]Ɛ[*w=,:^~H�G�A�gr����a*�űG�mZ�g~\��^��\�H,��4~e�w���rqȺ�Ե�ޱ��R�F�`��ɦ��-`�㭅����3�t��|��}B-t���G�I7p��
Vm9V��iaI��?� ͋���g��_5�����cn�1u?�����ňk��E���q���;@�e<S�_��O�Hh�U�ڔy:m�@/V�ߖ]�O����RD탣n$�J�Ԉ�u�J�YW	���=��6��Q��̈���e���\��=P��[c19���*��z҂� �:�m�ҧ�v, ���*�2�q]@:�va�F�K
��E|V��~-��F��i�ࡪ�x0R��ߊD�Ws�`�F�'T��|���������9�r��_�T�~����q,Q,r9G�����w��I>�G6���K�wGD2X].��ĳY����Xۜ���f�z��K��������!(?|S��x����oTR�"��~�,�߆�Y�{_�l��07��CQ֜�ќ3v[n8⫆d)W��1�m~n��;�������X�]@��8���m�{���x
!�|Z7zHsQe����o�14勃T�����F+Xح�v��>����Ԥ�"���c�i\�-�����y���ZIM�
�������_�UEG��	���Dڥc����3W��F Q�)nS�G�/���e"��m�tj�c`ﾮ-�~��%1�m
��o���r25�'y��9�~�S��\�$�KE� Rlc|��{S�Ŏ1�lًjĤ��X�ъ���N���1�]J8C����G)�=����ym���Q�0+��lϧ�+����9�Ɂ"Z=Y��8QpLR%����p����6�|��s��Y�������kr��L�Lrr+G߰��߽CB�2�W�/����_?����o����^�I0L)Zcuw�X|�?U����x�0j!-ꤐ��BOc����\~8��h)����~�_��&h;�b2�F^">�^&�,3XW�����,�+ݳ���ʺJ)�'����e�{z����C����P���t/K���Q��������~�:��
U寪��^E��c��4�l�P�;Xgs�����ְ�\�&?/�t��I`�t;>f���s4�cz3Br%wЬ������QV2c�$T�$�����NםCKM��x��ȫ�Mޫn����Rm���n�<�:X�@���/�L���r���Dkd\�hT�FB�p����"s�6 Z����}3Y��R��j�<Qـ�������ρxڨy�W�C�>+�E(l�\-��"�D"��k�Ir/�+E��}�	"3��M_�7P�ݔ1�	��	&Cz�߾$P��^�62z���xȵ��/D ͧo�d}�d�4�uyV>z&v�%3��:!��t�l͔ä���Td�sR)G�l[W���bF]:��O���Ў�L� 0Q��2�6ti���D �q�ُ.�������(�����Ŷ�XZ�L��aX�z�|AV㩲�4w�q�@��ƭ�l��¥}'��~��i���D'���A֟�i>��l��<��U��[��cK� �,�1؉;O��r���+�����0!�lOƇ���F�R���d�k�T?���jIEK���OC�a8�H�
6S���]�b(x[-Hx���Zl9�������D��t����-����ZjQ5͏�U�zjuOUr\i��1�H����U��/	��	u��ʿ��݅#��f{�J��dY����J ~qËuFT�.f4#K����C<t|,�� ������7� �h|��7|�q5>��%~��IX��j��e3��6#��0��+�2�`)��i���l��i���GL�Z��cV7�~.�!k\�B�X�4�����S�4����
D]�"Zfm������zڲ�4s?��L��9R*��=\+�{o�͍��NԈp���Á����4�rk:@�/�m�1+�8@Z�J���%:]��m��u%ݹ:�f�J���P,�g��w�����?��/8��
$��/�ВC*s�vI}ޯr��m)���J��w�a�e}.��=�?���(ܗL�4�� VZ���y�+oLH �76� y�jqzv6�?�e�y���"��ӂ4��ܭ��uɛeR�����ʅ�c�}T#{پ���'� Ӟ���H�)�T�}��B8��)�e�B�5�v��/�U48ca�6�ue����l��_N����F�n9d�t�K \�-8�:��lܤ��!c�G���p#�Un9���&�A
����j=�������� ���9�F�$����g�б)�}�]���(��7�m�^�p3ت����:�Q����3��Ǭ�r	8̒�J��dpfSV�ҲJv����/f�3^Y�rq2� 9�)��εÁj��ͨF�X�D�xg�x�^Ѣ!*5P���&��f�8A��JSȟc���h��y�*v~E+y�o�Nz�����z����QVg*�7��]�Ku��
��	giii�k��iv��7_"d�9Kq�+��Q<Ԟ�}]
Y'm`�S�X�llLj?&��lq!�%ߡv�F�ū��7�6����66��p�z�Wd�⺸�_�c�2F�61���C�����\��ѯ1pCg���q��]Lx�b�׊��y�RDR/qa��NI��]H# PV^k�7���Bb��,���t�����2Q�|}��Q�����5&���$j��R��4�x�h���.�^�"ۙ����DJ�?K��&>������7�,ٓ�h\Q9��"��b�&�i���|���)��<*esL?b��t�����M��t7�س�D]R"%^$�����u$[泐1w9���YcJJJZ��X�.��n���C�S*
J���᫩��I�u�U�����Wڢ;�����DX/�Fk�rat��n�g�z/��{�~�t�*>��NFf�"�.�����B�\�jZ�1l�#냳oT�_t��ĥ��j?� �vM^_���`�u�	E�H��n���u�i�=���X�0��E��9k�}���i�h�*?�3�#������s�L��x�N��U�<�>C(��U�eV�e3X�[a��O�b�Ⱥ��l��}h�q���l�����D��W�S
T���GվsS��]��+Qn��/�<�p�5�Y=�g
E��sM� ���vm�h0�)Zs�t\N��5�@��K_���kV��_�w{����X�}ץc���7V��cV�b7��2?���,����Wc(��*6�j��^5���C���6`�[����=`� |�	��z�D�}c�6�����ٖTLt�����]��<��Cm�Ƚ��ݟ�,��RL��b�doTc�C�i� J����b�(G(_-�p)���͑t#A�ߓ�W���s�Ϲ5�6�޺�E�����dm|{��E�U�.+��&4�3�\ �f�	����Ⱥ"O�P�%�:D��,u_����E��e�|��2Y�
]G)�7#�H�+�>k�= B�-�����gU��շ�BFm��kױ!`af�wsy�����9�poL(��K2��lݪ�c��M� I���؛Sꥇ���$��
�}��q��움]�b5�,Vd��O��)||%###^$w��;*v��cT=�(�4>P��hP�P�m[��h��Jv�>g����[��tq�Zi&���c�W-�iR���
�$ҽÖ��]�b�
�
�,������5(>OMAD��-�ck��qt�Z<��f��������.��O��By��8�A"�6�:)�?��w�>���wz��z�O������~"�d�J�u.��������'թ�n��谏`�qJw3���_�A��I�>�~�mBCH�ɽYEP�,Tr���]ѐI��>��7�ma��%�����<�d�z�_!lT��Sseh��͒��,l�h66>q�$V�f[�� o�nGm/qQ������]�tw�����
?�V�<��� ɕ����@/c^�q������P��t���z�k6W��9�?�oovC�CGϐ�Y�7�(�z�hL�W�h��&qy���=����=����>�6�,��_?Md���#Z!�S!����5�Nf˟�G��q�Ad�x�
>|�>���@/��o��/v��6��I��^��m�-��ԈVm�	q;Sn�o�e���K���d���4�X�~��#���)���]��#� �ˎ�8�Rko�9�W	�b���i�\cΓ����KY��~�N�D���c3��H���41k��y��P��NZ�r���!��m&×N�2��J����Dm����B�m)1�o/����3�^[��Ϩ�?$��?w��m̕@j��΂s�f��{k�U��n�M��y٪��X^�F,��'̸�0E�AW�~[�˱�LdM}�����5b�O6z �AJ7�V<nVS��5���K���������n���w��M~�|�o�˳&u������ժFX�@v*� �|δ2��Pwl@��X��y}�j�(�_F����+�$�
)���P��E���� �)د	^f��(d�zp���a"sJZ�;H@������%q� ^��~T�̴k��)�t+�uI��5A����smΨx=�Rl�(D�� :�1jU䡴��0I�
ko���Zu�<"�L%?xV9�z���7��B;�܋�P'I��جZ�����UZC�uEͨr�����Χ6���mkc���^A���c���6�sRo�=��mE^�HT�4\���͠@�G�?�ޢ���oV3p�����L�&dKK��aI��P��R���Y\d�Y+�W��D��LF��hy�`� {W����wq��1�%@sp`��黛�2��[��UwSpu2�s��.��/�9�,)yy��S�m���W���/��.�SZ)%��~P,�[G����d�5���!�ߍ����?�V+�_^�i'��y��Y�6��?�ߥJ �+�� �3�Yorp�!Ⴢb`��4纾�e�*/%K�kҏվ���ZӽY���O"�"o�F�9��B
�;��_Wԛ-�)�?���$RZ�.�n�4򷌌�,'w��B�E�/���/�B8��bͨO��H����$���(#>oln��Xw7�2�A�{�){�����5�2���gCnN��K������ ��� �3��h�u�*�Bdy̟�1�&����8[2"���`�稦����|b�f�²�ⶤj��i��j�ÙN��_:<f)��|PPЁ��L?i�׻�w�Dg(��fި�Y�?xT&��*x����fi��2�^?�
u�����0�_A�F]�q8��#E(lg)�����v��Ry��M�g���Ǔ��c���H���UPQ�B�u��0��ݎ ������dV)��;eQ^�S)|�g���[&Fk��u��us�ß��8O��b��D�]޽sx���o�Ҙ���j���2��/�-�ٿ����s$<�H����i�!����Ki�\ 
��}i�Ł%�@���Ë$�ۯ�����O7��L��*zw�O����ס��'q4D���$1ā����S�uj��s9F���Q?�g����+��}=Z�[MA*��WN$��0�Bm8�ex��P���W��ۖ^.0����<���X��g�Մ{SƆ�n�Z)�=a�c���Y������R���lh۠�:���[�ڃ�C*�i�!a�Fłr]�A%���R��oVX��x��/�>Y#/��~0�4�H_C���7�:����ٝ�$d!��..ˑ؛䁥��=<{��]��׫a��-�����>�o6s�5ro㬟�G��T�R���*K��G
J�h�;1Đ������"l���9�V������F�B�� Z-vG^������yI���7�GZ�Mx�7;���q
��I�+�`�P,L��J�4f(�?���b&���;.3���Ѯ��W��@φ����pg'�!}��m��ߍf`ApЕR\[X���mӝ���̈́_�n��@*���j�T��DK�!wk[�3:`���Jʮe�N${�p{dmg�q!�q��m�șo�!0J(�vx)3���4������[��l
.顨6���.1!�7I�V��R��8�9�_��M_jjͷ��?��3����{oѓH-z���#A���E�DD���^G�ޢ������{}g�������>g���>{��hM}�nY�0酜�� ��Q��������eK����6��G���	���K
���Q��#���Ir�'�7��?+��`C��c*�}���ԟxz� v4g�KE�&���k��q���UW��q�{���_�ld���w�%2�p�S�>��{X�xA:Mڛ���2V\�]�ꖕ�{0	<1y��o�yz������	Q���6F��r}����u�8Ib���b��م�����9�Y��0_>�鿪��*h}��lh��
v՝���{�a�حƃ�J��8lsL� �A�W�H�8�LM(�F���$�����J�`MQhN*�����ɉkso��RS_/��9ѹ+w���5�����K񼽪�C���_��_��[�P�e'�e�餳�f�����LD{�\o������Ǉ����V3��Z�H�o�>��ײQ!ڶA)<` �ŏ��ɶ��e.�����ן���D���IvK֋��p�ɑ�x)A�/�Zin���m�'ci2����S<��ñ���z��MS>�#q���#ҝEz�p��[���y�r�`�"/dL�8�N���,����n/�t�ղc�/K��zP�����o%��:��x�j�%؍� �V�̠a"��;��K]T7�Aᦱ�;b������P������dY'-L�w�@[:&�����&%��+�V�fZ�'�?�J�z��ٳrM��[���){�Lju|/����K�3\���Nd����R��|�1
��a"�z׀�J ��Ճs"K`m�2���G}���_�䴡ɔX7�*����������������h\����qR �)�/�p�|;r�o��tص�e�ӱɃ����֛�}S���JFi����w�����<?M���-�X�H&]�b棉�.��͐�>���Z.�)�VU�z�N����$�MA��bykC�!���@xN!��E���f�9���4�҂z�rJK����1������;H�e|��&�/�E�ȏ��:��ೳO�<i��ߨ����ӣ<::z]C�C�TPP�<ۥ/.)Y�9;;yw{u�,�E�,���J���#x9R�UY�R�&A�����&<{Ϧ��~G�4�:��J(��ۡi]����0�_Z������|�_��;W�6-���x,�8�8�T����w١׫m915�o2��5o(��F!'%�˼4�A��9�h�q�3^��)횭pt�턲�ؘ�D�����ls��QNlu���!��$D ��k������ ���6ʒ...����[��=N--�Q*3y�� ^���Da!���(ZR�y~͉z�?\@(~���^�fg'��{/TBb�	+�B�*Vf�p?4�ef`�w� ����n�g�ms��g=J�sx|�GDJ����ʿ�ޚ��-���8���%3[�ɯ종�����{$%$F����y���x����y�I��B5�_y/�F����`pBb������~O��^�/t��+�u�10D��奲��i�����^	�9�3$����hu8XW��S��j��X_s6E󇗻w�F�G���kdX���"'N&7�(�׸�n#�$>s�� ,;���|;@c
'٢����`s8s-��gr�3���^N�Bܾ���~L����k�:Ȼ�k�:C�*�Tɩ�6M�}�<ݍ�	�9����11�h���6�|��SMъ3.RM,�$,8rd�F]��6:@`q�b�����n)�*�8�6<�+Y�7u�7u��я�U���g}䎈�.Dsd�O7e��/ ��3����4��mz�m����߸�^������{ ��Zh�|K�u(ޗ˔�J�� E�$)�(��ǵ�Pg���ǿ4�����n��NHBW�=,��k�����Q��T~g����r5Vr#uKR��3?"N�ʶ+j�氧ɨ1*!>���x*>U��jgdW�}�����J�r}�,ٚaV#"j�{Je>{~<;1�jA��H�b.�<Uf�Fn`b�(���\);��2���6��K^K+�y�De4ۏ;V�|���8���9F�4���ϣ�	ƧD�>�*}��S+]3����~mu���ĕP��\�����󾤤���­NmzBB*���F�b�݁�ZZZ��E�s���?�v�B�b����7����yF�B��T����D�M^�	t)
�t�E�.
˰��+"nϾb�2����`�7��K�;S�!X�}����0\���u�{aZg�{tɸi���]�x�}c�wXi�����@c��ø�'C��*󋺃/ͺ�����5x{�	`�H�<id���7�pm���KeTB6
�#֡�6��;l�b���[��H�Jy����&��.���š��''W���> ��k���#~�q.�=̬�U�Q���[m�9��=��'~Y���[��k��D��*�^д�qՊ����e��
Z�3xun�2]i��������S�X��|�w�_��o	��a\�DX�X�%$�n��M�*M��.�ɷ��V���ř�ô.L"�F�	i����x�Z�1���V�m��떇�~r�
O�-I��!&��w�^��={g��=�������#��f���QVW~iB[�;����V-�kg�:靿UL%���AV<�P�_����rs[�a��G)�~����V ��mp�Lq
��ފ��v����N�w��K�t����U.���u~�wH����dSq����,5[=W�hM	�[�������mO � �Q_R�_�@�gs�w]��ԃf#�sw����J������f/15<�?�.&�uc}y�.�� ��NqI~��0�P�c����ٞ��2�S�G� h�AD̊�N�;`������mvC�$������g�˔����|L���D8w������;��b�diGH�N����*�\��K,ܴo:H�ј�^;3���6h��K�g
�C?��u�֨`cUz�jH/��W�oV��+q�A��*�s�tp�TQL#j2�D���̺VfD�B��k�<������W
 ~W�����.1I�T|���F<z�yMb���	�y~ն�C'��뫊�����s/���S����IB�]0�;[8q<��q�FGE��-� �ڽ��
�HL3酩aS]�Y�WߟvA~�6[QZ0�-EO�ƍ��s�c�T�"����s�uT�����)<��'BXm��6����f83.�	�Em`�j�h6�3�c�˭�����_F��/�z���vgy#�	˳ù�_�{�B��/����Y.ꤟe=�	28�=��貓��`�T� ��~��&JT˨`3H�}u�;��η��Q�E��@�zv>�4

S�NK~��Ws`�b���1��ҹ;(���#г�8�$�|�e�0y����&�*�|�'��G4�q��:�Vi=����I.7���/�qŶ	ևZib&����OV<A<w��)t��Y��[_���FD���yH8x}�4BDR�S";P�"n��;���G��X�!��(�:�3͕�(��o���&O'4`O� �;�^s8����uv$l�:�Ď��D�gy�v�����"رԅ�Y�W�i�`���1�����B��|�͟��|��FU�kjz'�^c]T����w�\���?�:�||����k\e
��}�(����T��뇽c�7V�վxϣUU�m�L�x���`Lpv���U_q 7�6b��W�����_<��	)��[�u�����п�-�������{1O��A^�����O�Ž=u��#��?��Q�Q��R�x&ɄZ:��+�Lsh��L�\Z�'��7���Ik|�U���)ڣ�ذ���f��$�^��i21g��Z'�#��������׀���>W�s�7km�A��ѡ�8R�O�D�o7�bv>bk&=A�|I��"�<�m �u&0�랡�o��nu����:�f�KZ��xEX���{��
Q��a�m����C�-�t;�e=EV��B��/Q�ᔐ��8^��g��Sşp^�މ��t�����R�bO�t�ssv��!	{�Z'Y����06jc�q;��.��Aeo����w�d��k���.�:�[�Cm�3�Q	}����-m2ch�n��߶��%�\��?F&~��L>|\�����f��[����3�+"�����(Z��_��Ŏ�	�=M1b�\�/^�(�u����R�2�YvnK�|+�g�T��n�B$��x��H&g����h% h`��D��ﶷNN,�"���`?-��N�b���y-�t�.,��s��}��H`�%����&��ٮ�3��?e�_��͒B< �}7�����; �g&qN	�b�G0��=m	��Y�������q֨�~ei�7bIE9k���'k�F�������P➳���Ew��HD��j&Kxx� ��2ݚ�8�/{��5#A�߰�y+]���y���I��3�}��/�l��F�� �$D�O~���W���J��%�&�?H��Ox���I7��,��+NɿJ� �#Kd�����D�����*j����d��rE��A��	�Z/�}��H0Z#P��3,>��7��DK����_r��,���9�d�L�p��X]_�J�i�ãP<�q\��s�~��S�m)\��Yij:�}rIPyDр�f�����S����{�2�S�$�NZ�Qڡg@@�"/�Ct]�d��t�V5�Gڜ)�i��Հ� Zw��n�z�����q*=3.P-��\���`��W=���,o}�`�6���������"*�_s'�t�2"�y:4�b6r�ik��Ͱ��S!�Ѐ��	�ah屵���Q�cQ���4���]G���!��	�\�%�Q���p�O�J��?/�'�-S�vuay9�*��6<҇�n���!	�d�������9w�&�wJO|Y�$�bw�a�(�y��H-�����|bp7s����@����*X���R{������Y~y6>zĚ Vǳ����F������Y�ɿ� =�(���Qg\�m��Q!+�xDb5v���x��^ ��J��&���j �jqK�fSƿ��yC3(�؁8�Jz6�̕et�_s;���"�7!�uT��C�!6�~�{1��j�H1�����[��;`탬7t?~�>�z8�aq�{u�7� �o�����Õ�f!T�Q��_�R$�<�*�u�z�W����/�N���)��z������Y��&���M��X��3�P�">��0e]�+���00�����M������6/ND�����B%��h��I�d��`��µw�C����s9��X5�B�Z����~7���?����6.`����_��"�1���n�6~�����\�Ĩ�&$�?�U�M����Nj��CAf)�%��r�z{��0��%��ׄt�2���I3.,,EJe56�P��At-��F��4�&gg<����Ʒ���²�EΧ�I��<� �(h�	��$k�sB�)�=$~#���0���7�9�/�q,+�c9��ʹ�U�.��/��E�S��0�P4wa���n��mFU�m�b�>9n�ց���ި�@a�����(�P�X�l9��JQ�B�2WJ&�������L�H�>�ϐ��]F-�9�{�ɾVR�?:>�w���s� ���r!�|:�aS����d��s�rR���S��I�Q_�L�yc�)M��i��n�6f#iqȘ��ܙ�bO_���2�����ȟy�8��V������s��fۤ^�|��Q_����*3�
۳��8���6#�Gl�Q��t�����ŧʋ�:�:�@\(��RS_�s�%+S0�+Z�B-�Z-�d�b���\#eggg%�o�[O�ߖ��&�LG��$A�G����P䯞mb���23GJ�*K�ﶟ2�l7���	qq7r�Q�[��mMz�~ �?�J���W[�"�X1rL��6%㰔V�n�����c3�=!V�����t�(��.�T�P����uض,�D��6�a,H2� �������vG7t�ƒ�M���ݙ���ȨH�5�v	ʝ0���zT7D�a�K��L�SpGQ>�D�eJ������ ��(�p��1e�9�>��b�N�N�z�N������I!�3c�/zb�<������V��VPٞ2�������b�����5�k����@d_<���N��^GlƿvHRB���#E�Nr��:E	�$�ϟsw�iDO�kp�A�L��±�'W敮����֘�=��;���jHNN-�d���D.�j<e`B�8��ۡ<g����>�/���V�a�q�
��}����FF��O���A�^T��{��Xg�'��#Z�}+��|E�m7�ݧVkE(�YG�2S���'7�SC�.S��j%��^�u�[��<��;MJ��A��rr["�Q�u&	 ��G�;��|�;'���s��Ѥ�E��D�����Y��؏�w��O��o����g�G�֢m�D����W(x=���o�e�JӊǙ�������A+}_s�4G�ʁ��D��OH�JɋBŐ����M�x3{��*��}ʇ�b]36�Y�D�C稼OTm�-\]u�
9J1ҞK�����=��l�����ޟk��O��G�}b21�#d��Ɵ�R����KO�o
������Q�m-�����M9/��l�|:P��ނ��݃?<��q�VB�RPT|��>���~۟u <�"����ayE�n��2�G�~�7U�^b��p�s����xr�E�sw8	�����?��ԉ���_F1�����T^ؙNT����^���:�j�p�l*A��o���;pK��("�ݍ�w��i?x3��F4brfU���0�1�ƈ�o�ؒ�� �*Ҭ�b*��Rp�03{�k0={z���%WA󆳺��톂��L�����Ǭ�h�i�Cj�H�M�fǩ��$�t�l�lϐ��ypu�=��d$�ӱ������5�x��Z�4���8���4���AZ��dlޯ�%���Վ%{��&R?��U��o���x�B�)�@(8~T��
����'+}�P��� �AVzZ(�,���_�A!Yx*A��]��d%̹SvOP�[��A�x��k�O�)���@�pLL���LS�u���W�6��im���������G��C &��9���YE}/]�o.$BAj4E�y�Q	�6�2U7-�a�sk�2R��P��fIYV���EW ����wzQЛ�����6����i�䯏��&�D��֩'d��
ˣ�F�P�#W�Zɦ���'Ϗ��y��rG�@0^"RR�XN]ug;����-�.:E��'x6��Bg���{P	����V�y���=���]�k�~�i���Aibrk'��1:n&ߧ��YS�):ByYg�҇�?[=l�A��"�5���!0k
�{�����o��H�[qiq������ɷɩBڃ!������.�.���R�u�X���
�:�f�ĢQl
�� ��Q:��\��[	H�Z�����}	��趤|�P<!�/R+$G�czT�j�>JIύ�B����@�dI�.�ܦ�&���xkC1rw߽]-���]�4Aġ܊��|Yv�0����y֩NX��b*�`��<�x��	��>~�ɧB����$,*�r�܉����ú��ۗ8��O�ASL��s����Z}1k�F���t�ǿw�~KD��t���,nU�[-�c�Iԕ���G�|w7��I�+J���i#�&��5JH�5s��?4���nJQt��uqq����9�T��Nf��C��Ӳ?r/D>�V-�E�Ț%��d�N�3�C�� A��~��yFp�A��9��>f�,kEC.^xA����S�ݩ�&�0�i{�r\�x���ZX���) ��Y�!<�1=	A�s������^)f��u�Y2�K�p��Z�bl�������gB-�sr����!Q{Я^��ޫ?�P�L�'�[;�v��1>P�ѣl��л��Q�αv`���&���7؉���˱�{¶L=�r���zG�ϟ??�?W78��7�<�$����	�gY�\�qss�]ិW�Z��C�E앒��������F�ɣ/����,أ�G��t�Q� ��9i
V���\����C1��A^�k�$s�	QN���,n�Aq"ߖOEc� �k�1w'�@�
ӓ��d� �x�A<��mu=Z��ˈ�A�����:uvO��B��hZ?�:ԝ����m�Bg��;�}̄ǒ�Y{p�S�W6��:���N����4�ߢ>[���QbX�45�KXOZr;M���.U(.VT��K.�z�/t�0�`�@mO$����i�P]Z%��YM����6vQ�te�[e��)!�j+��O��gE��uII��]�/f�=]���9%!&�@9�Z�\͉>��*J!J�za����m(]�r���2B(yG?��c���6V^H��GBˤ(��yp����J���h�/��K�
Ry�!�5�Pv�tb>�R�O�YP��+�qm�,�!��Q�ns��/��I�:��K�n����;�O��~��7�̞m�B,A��"�}GPIU����8�@x^�o!�M�2���2r&&���('���Ŷ��R��'$t2��n����Q�8�i5��B9�)�i��@��(���+7���h�y\JHNOO�@�iT���9�`�\�\�/jӡo("��~�����k��2�����;�o��^?��8�A1�� �hv���w�vr��L��أr��_Rf)Tfv��"����]aP|������@ ��>���y�6��q�5E����[J��z0����o�z��H�/k�cG�P*�cN�p���ÏF�2{�0���5*����z���x��8!�O����xpᅻ&���3...J ϲ���>O�16xB8F�lO{��;$���o�#f�����ΨSk���.��Oz,R����������n�u�;�y����(3�-,@�bY�؏陙{ �:iF_�
��kQ&�E �X�ޛ�n�3�<�IR��"f�i�^���}�V��_��e�(�ZJ�	}Fʕ(�ѥ]�q���A�Z
���˸��QZ'Պ����7*�����l
. #�CAx���H���}�`W]�G�����O�
���ԝK����ҹ&��� �NO�'^�}��x4Y�n�B�syP����ҌVηF�=�q��ۛ�ڦ8�ߛ����l��_tL�F�L2��_n�����5?��`������4C��E-��y���l�껐u@�zt�r�O�b��F�i���Y� �����F�3-7{Z�����\	f���U��pv�_|,
�y�g�<�B~O���q����uH%x���\�Ȧ���*�ל�ڐ��Lby��U������k >%'o4"onz`�n5[;_�n^�0�L�uyyt�8���ߛ�����=IpR�j�K�(�ʮ������!25��R򍅩���h�>d����1i5R&�ht����7��7l�ZG�'�S���pjg,%h�8ǰ��6+	������ag����V�9;p�Y��Ly��,�����ݓ����,�Y�#�a`d<<ZS��	��P6�nL�e�e}L�>#�Û���p3G~G���Q�*6��+0�2(�D3�i����F�0�<k��<y�,�$� �X�呣�j�#�"���ޫ_j�T���K_�#p/6�ŻM �{n�݁{X#$����?�ﱏ^9:�Ⱥ+��r?��OD�ٟ������=��I��8dؖ�ާ?<7���>K]
�۝���z��7Ω�f�2�\{]��YK�c�� ��i���A¶y>L�ub�%�M�1VQnh��.Щ�DW������R��g&��-���>�z��5K$����qa���FIF�����j�_�<Jc��,�aN/���p���1��E��~O�a\3hO��D*��J�[��t6���>��L��V���p֚��Q���g��lR������X���]�m-����c�j�3���lw&x��nP����I���Ѫ�?�����_�u���k;�(%Y�����sbs�7r8Q���t ��P��B�զ���c<t���PҪ�ož�*,N����)����n��`�A�*���%)���3�)*KVr�E�h��W�\�=bz�h㽥��!HK��3���%��@)
1�u�wWz[E
X�L���8�&Ys#�1%uT���Z�˞��-G�5��|�5+�k�7�=#O�V�5«+_+�Szn����t�$WnG�<��Ep��V��D�;�T������7�3��U��J�C;ִ�/B��{@�����ܢ�vL���0�S���u�^�%}h@i�Tpy�S(
���$������
E�Ũ/��<- SR����f�qK)j/����/�T��Y���+*#�0��C��0e}ߴWs4u�(�s�&��B���Ɗ�єV;s��ot]l��(f�����z_m�-T�3]e���B�B�,�	7j�@��̀3**.����@��`d����� ����2.�Mǰ���>��6(�=�1Y�5!y:;�O>8�P~K������k��Q��@v����T��9���^%�z�-��4xY%��:� ��c<��ᑛ46��!c�;*�V���[��J���7>��ދ�ܿ��2w���h���u��7EGfS�IU�,���	u�t��?[8��<�b�zs���Z��p?~Y�jc#37/s�&ݘK�����ڴ"OZ<���C��q%�6x§s���5���{�
+��qI'�凞TVLD�'"b�nGF���g���\(�1X�Q�p�����,hS(���u�Л�P�*���[Z�hm}�CU@��-�^�Dڮ��ݓȋl��ǘreؤ"@���Y�r�������gi����.�(����}�G03����S��A���)t}�#��\��N}$����qd��5sz\[�����K	���Y�~�dU3b^G�� ���{?^]W�X�3���x����b@�;�k��J��&d@+F��$�#���&�C���� _�@�0u��8"P��ٷ�?���'�*�#`#��L&��	�ΪA6J�9� H�ğX��2���MYږvO$B�Y�'2�.C�;��Q:Uܣ���?pFm�d�h��ɗ��\���X�o�����p�!"��&Xwn�����&˹�Y%�0�`��)G9!X�h��C�[���_L�R�,�Гף��n}S'I��(�D�P�e�M[��]�e��:�5�����`R%D�cgVN�������Y{-pr��<�WC��sd?2�E���H�l�'���w�����c��:��^��fӺ1����y���p-9ߔd���D�z5�7�jQ&//V▩Ǧf��|U��9��Ƚ4`�ӗ�b����[o�S�������M����-s�[,WX����$��1\�!sz?��\�؅�Q�ϟw��"S���[
��u�9f��<g�8	��8r��r�ݖm�D����J�,b��%�+�v�8_Ё�}ű�ߓ���Н��Z�N��h�"*0:���ھ@�!�7�$;�:ǅ�H|c$�����r\����?��A���4N�E�&}nh�V7�>f���Z�̗L��� �C� 
�芧�FȪ�X�����c���'>���~��4~����M�X����#	p�c3õ���w���p%#Ƕ"7M�ьR������͐��x��j�]h}*��a4����l��P�}	�U/[����xS���12}��_�=��d��˧����1[�l.�5^+}�2�Q;�Ȅ��vl����:��׿�w�qϨ�z����ͪ�,�������;���X~K���T�R"l�_�OÓ�o�L���m_��9��b�v\�L�5�ҩ(� A�a���FU�{����\��O�N�=��p4&t�kK��N�%��Z!B��&VP�����tx��"�,��|���ʼ�m]�+��7�:�@�����C���u�oR��PvOZ����+� ��(��F���"U
� 8�)8/w� n��:lZ��	��VwJ�Mu��tY�mf�o���"�:I5]?�p-���H�E��g���eyK;S�w�x�SN�����^9���~���Go��A���b�����>zm����I0Y ���冿�H2%���M*�Ŏ���G����(�lOk���?`��"fu�8\�E��w?��t��c,�}w��A`�&1�&���\�~�G�r/����H�4!f t�4�H˒R��}@&q����ݎ�.�C�<f�ߕ])���(|1�	�1�$���8��2mq�s�}S��5F�J����V �U��m�����?��~oetmm������� �60��I�9'Z`\`����{κ"��{~���[��N�S��[ y����yI��U��!stK�����#)���Y�$��)�(.� ���%��*dF�\���2��'Ŧ��o�޿�0���!H-&��dڋ��Z]���`$J��_8��22�tiL�T|��_�_������ݥ��7�,n�o�Ϣ�� c�� ���ȸ�����'䖎�+Wq�A��}씰��?T�%^V�E���Vi8�w���ʠ${����]� �Tq-k��6{��1Kf(o���jOk�aaM��Hy͛m%���T�7�Ӻ�[pGa�����b�8G���}�o��XX�|�ú�+c�+�Bfy�>��N1��5O�,e<�%��hn��^7]�8z��x�2� [���x���T���oy.�K�|y4������Ϙ�.��]b-W�S� %]�do�g9V�{����N1�����Q2|e��3o������%� �7BXs	s~D�vy`��^���إ�Ҳ�e��ܘ3�{F�>���/��>=Yߜ%y����%=��Z �ƌ�=&����I�ܽ4����[����(��#'N3ÖK��ѣ���r��?�!���O��3�6̘2"�Cep��/�I	x�qvGv&�����K�犜��Z�� A�����^R析��t2�l��]�f�݇W���Y�{z���*�>YA�jΏ�~�V�o�lk5ӸO@�m�&���~k��g��/��f�SU�[aC=�~�o�'����k_��,�0UiҞv�o
�%e{�-b���W�k9E0��l7�9H���E�o��dR7�Z�@��9����w���(�&)�ft��P�����'���Fe�N�<i������1l��*D��MM��W�,�Nx33^d�4 ��[�6l[�l���ħdsqL��w~���f����'Wo��苆Z�N�&��,���$PH��^��ͻ�<���Ր���/#�R�0#����X�G9�ԫW�m�ug�4r0C�y[O��F4����4�9s�%�,����2Vh��I�t�����:�A���[_q�y����Gd:w?yG� >gA�d��v�Cw��! G�	<'U��:J�/Ѓ&)q�Ò�l|Y��mV6��T���~���yt��y������
	E�`└��Sb�FS-��T0g�M`���c�c��&���v�w.��,����b���̴�.�Ż<�_��S�`�?�C��k.A��Ϟ��
��B	��cIᘙ-��.��Zy	¹�f$����}�=��e��[����Ãe��÷UUU�����7���!242J��lq�hn�Ӻ���ly�`�9�?�a����y��筨�����"��b�����90�����J��[�7��������[1������y��@Rn�*��0�(|�z�/�i��LE�&�h_m�O�>:j�h6W�3=3}{Gǃ��Tn\�Sޤ����u����9����u�9|�|qd�|4�Z�!��z�[�=�y�kr�[���]ћT�?ۆ�����;��B���5��JI �d�
�=�7m�C&�!����＼�g>�揿�I$5Rb�/�y�����u���'o�!�n��q�|A�r��	o_�☲`n�880{[�'�o)+#��<��o�_�Ei	G;���n��}_i��q%x������ԃ��_v�x|y���G��K��Y�V$�f|�[��Q�u����v��ʔ�Ge����_�DCK���c��ż$���jlj�éc��H}���Я�׫����{����o=��yX��X(��{]\[]<F�w������SG����F*6�܋��[�~8CC/*QLW��m_aʥx�o�Bg!x����"?�����SR�H�oRgG������K����,�e��/*���;L����F����ˑ%���)K�<*���R�o�>��j��lo�V���Io��IYt�xp%f�ڴ '{#�%�"d��#JE-�5Jv܇\C�8y� ������D$�9y-��|J�����D�OG$E��n.�J���VzY��67mm5��6��SS;GG�&���]��.���1P� ����K%5�P�g���yg��QW'RS_o����R^Z�ty�1��Z�x�)�@��P������.��8A9 ����wB3�xg���A�|ځ �p��W���Ʊr��֮�Q�瞔�5�ߚ&�h9�!�E=P���vg�~_8]~�3�Ǽ23Q�y���n�!�ڧ1���y����$:&&�=C#�{���
�&�6�_G��>&l�M����{�p5=����v�j��z�[�g�&��Q�wr�(���aPe�����b�%܋!�T�KQO�0G�Ƥ�`���^v�Q��;G.C�c�y_��na��3<=g{�������TS=�444j�k"��PY�B�¬�p�����:��{�T9���p�o&-_?
�O��֖�I��k����o��˟��1?-H��1�ܷ�ߍ�2N����l��^��������%$V[DSK�d����|���"έI�9�?��Ӣ�iZ��W�E4�?+��'p3�y�[4�N�����»0J�j*����ɔ�O��{�z�I.T_Gcch�e�Z:7�v 5q�MGs#Ύ��DWـ�_eA5�z�7�f����Wv�%�8�(
�ׂ���t#�v4|}��(?(p���XA�-���>8]��ޜ�����>kY|M��m�<m��#m$���4�{�,^Y�̔��eE�sg��p�ͯ���{�����V#�sI7��7,�S'���Lہ΋��4��_e+/���H��_]�t�9�K�<g?+%|��\����Ua`1<ʯ
p0��9ğ�y�;��ʩO�*tǛ<88辣�8��;X�L4v��z��n��q�~v�K»i�C���$Zv�RS��P{rޏ]Yڿ[_D������'���[H�D��Q���G}���es����=z����676��2�fAߞ~�;�����!11ۼ��{�G������ȑ������:G�h㤠�!C�N6��W�^d|��֎���r{�//�܁555��ՁD��0�
���P��H
G��pi�pm��m�Rs�-��#QQ�bi��0�g������v���}�⠼�L��Y�-)�́��X�:N��ꣾe���*@�Q�'	�t)y:m�Zdü	m;�J)�b��U��g�jȪ��*��)W���-���?ƅ�� #Ejs�gz��j�����6�2��.���|�����G�B�p3�˭7�|��������//-$��`�"�u��|�)�n�,�]ˍ���G�PG�9�,��X;&���|݌�<ވ���2����ν��0L�R�2OW#& �ss���j`oَ��/��e��_:[��.��i%�z����������-��n����{\�ܭx��˸�G�ߪ�5�T���gf�����#c�Zh��z��S��keg׏v�U���]1%����>0W�ӗ�s���`5�j�*9�Ih)��^�[��|RdZG@���	��j��ׇ`���5&g~��^��[��u��X+��6�.D`�j�NlM4��6����H�O��P4�I0�+�a�.)TX�{22E���ھ�8��,sNJoI�,�W�|�w>� o}�X��i�Wo�+|i��H��k��5����!�<?�0��ͧr0 �d�e�06��	w:0@EM5�������|:p<��〮2�09������4 �[��B��P��V�ǝ���@��]�紿��|fKۓ%E���J�|oFH^35P ��=�iqC�H�G����ސ�VJ�;�l
v�8?(	��k^��<���s�,U;���8����S����HZ�?k'I<��檅��~OzoN���
��%I��3h�qO]:|ll�B2��H�����fpa#��w�y���"9)��&�4%+,��x�t�lxU�ҹi�8���	җ#��C��Ȣ���]n`z(��?�mo�	ò�£*�	�P�+!DVU̓�����'a�$�±����"�bn�L���y����_�.�u�e��ޓyΆԅC�_��M)$��h���u^�!.��!0qM���LF�0�� �TS�)�z�sű5�Y�D�{�����F�k'�i�X���_��xć 6��rź/2�#m��쮞�a�!!}ǡ��M��ݪ�-��TH��Z��;�P+؈_���䶋�8Q��#�8QQ��ُ΁?a	b5�_��e	H6.��?u�ם#�Sp:n��u
�yo�ݻ����*8��E)HP������)�-����+�q��"��ri�����M&�ZC}vQһ��e�?�����S�Y�w�O|������?BN�O�Q��¹�$]Jٵ�f�/˥�����9��+s֕g���G�u�C���J([ȦP���EHFF8;��l���PvI%�y�93�Ȏㆽ��-�������p���y������~�^�.0�7��N7�t�TE����8��?�Yp��ޝ����~�IL��'���wg�ݛ/�Th܃邟�"}<��N��Ê_�M�b�H��\��m$Dw&N�>���t!�7Bk��G�]s�zo����DQw��D;tO�+�5$T�A��/�ۏw;���
�{n�k�.���!<b�m�584� �c9�) '�l���
K�����<*�k{<㩙c&X7@[N�8%w�5n���vi0���:�����C���oF��I�S�3=��{�+j�=��OD����t90���qp+m�X~��lA"���:�y��ݙ�!�sF��_*u{8��gu�*]W� aY�7|V�u�"�S7��CL���^�Q�O�>���,�~�'ާ��dgm�3�+�fVV�}.���O�);YӉ'ȿɀ3�;�wr�md	�̷cy$6���(��~oj�&���Ϙ8���|��.)kOK�m]�$KH2�Һ�nv.���i#���%��fb����srU$�i�R3o��~!��7���P�K�y�d��U�:zs���~���/R��v���:�X�A2�B�ٹ 2]">6��ٌ&bd|+W%�Jbbbq�˳ Kl@�T�{
�%ꅆ�Ʒ�P���_��`�*b�[?���(EQ1qm��[���R*�a-�~���<[&3qa�q�9H��m������s���;V �N��fu=��=o��3��%����1�ئh��LȊ�VB�b��I5�:�${(�*�{�ݫ��N$θ�q��+S�@���n�㌑Q�������j�/Z@��|.1,���.����-�y�F�3�H�����������mCE����dM�yܴ��7���Z�]�D<?��M��Z����e�JN�u��>6��(�ǻ��6ҊJ���Uq�g��oS���bb$��Q�]Vv��^OZJ*�7KB^bb8��}�e�3����ܣˑg^���SԤ39{��ki�o�_9B�B��8^>�j3淍2n�{����N��������m�Ý��t ���>�QB����_׆���SWpo^x�d�5fl� �"����#�̞_zd���&�;�Ւ�j@^ �9���ύ׀Y���"����򮠠�$������YV���W+�R����_��TUk>{�K�3z�U0�`�ڧ��6�f~�a�˾A$�W)��\T=������U���'�jc'L���]7V�A���}� ��%ր����`!V�h[���_�dq���Fɜ���z�r'��B�R�4�>�
��W3�1p#?�\W���rX��8h���P&�?��^K�����~�K?�7h|����D�nd�8��?e�cOR0#��2�����k�B�+�G{�uc���CJJI��	������������Z��>x�e�Qڕ��g�SOa��X6J���;����K,�9<���ҍ�߈b�x�������'(��ƷŁD���������T�mD��>){[�L����������w��{��&�F�/��R�;ż�iu�k�&����߉%;�w�siǮ�^�}Y��޹�}K+\��T2J ��IsU0ݴ9}v���e�fO����T��3+��Q=��X�0�2��5.� 6��Y�ҸM��q+� 7�*o�T���<Q�+�;e����`��?u��?L0�v�ػI��b�zy�dqu��C�%�.��>�/	=~'�T�6x[ǐKB�KU��Sv����[�q)�nzo����K|��m�8����R�`�̔��:` 1��I� V>�P�ȥ���:�| �d���Q1Z�2�u�2T�,99�,�-��l`��t*�"���t��~r���V��D���?Y2�:�^3��q��aQ]�I�Uy�?�F�{q���wl-�_s>:��V�_u����ڗ�0-�gϤ�u\&�(q87���R�H�rv~dd�?D�WJ�D�I~��΂�O� h�>�T�$uU�6�x�	/���� G-U��$�R~��z����<e����򹌆�
Z�'�n7�b5޿x�ٰS�@@��&m(AH�r [�{�� �3�9E!����B�E�_�1�wޑ���Β+r�8��`}tR7��͐v���`�o��Ԁ��t���G����tRi�8�#�(����t��ژ�J��')��.���:�
qzwy!q9z?o��C���O��'������D9�������>�����r�����T��Df�G:���s鹒ᱺ̱�Ci.���=H����xT^4�����,s..���-�k[%7�Vs��џ��L��ߕ�� �������t����6��HN��T��$�V�v�]o�ǡEX�#�R�]/0��GKMET�CV8�^�)|���|X��^�����xA��~G֣D�&� �.p��t	_�f؂��WVA�^���Є+�K�ܖU�i;^ի�1QSS_��P���#^��
e�_�jh�W0������l�z�`�h,+N'QV���V���';�n0����l
��~�f��V�#+r��3i�g��m�_�?L(��T�`�]t�j|/K�����z����r�Y���eF��f�l�gJ(����6�;;'gs��[�W;	4.�[7D�6�|���X����8zI�AȐ^���qo�N#���ys�ٞ�MT�퓿�x�C�xi@��ôz޽����ф��Q�X�Yէ�<J����F�?�����*�����j��W����Qɏj@O�p�
�	�\}1f��Q8�Q�r��ǩ���דy�)o�C�-�3�u��A�U��ؑRWO�e����č_�>��M�Pz�-w���ޕR��N�Z����Q�^�x�Xkֵ�|�]ҭ���,;/(y�+��������,������(�N��6�6�_��ɏY�eNI{���ֹ�+�(��y"l*l�"W5���$�fy�s��[��m�}��xA�����x¼��唶l��k�׹?;���+T����N>5��%���)O�l��g;F��5�x�u����[݋F�ͺ�	�T
�D˲m��uu_�wn&�QG�˅Gu�\�q���b���M���j'1��܁�YK��ҩ��'a�^��^G3.����������r��������A���2���eWq3F�/j@�V�����!�Q�^�����9	XA���QO?�-����X��bZ���U-��r�?.��{�=]f�)���sn^��k۫EGr&���M��<6l�4��kW)3+���ڇ��4�r�6��b��}� �;lY�yݻ���<�^T��^TkVҝG9:!bVL�?��V�-��K��v�`�ԍ��ŉ7)��}6i�J�@>�]5��c4�ː5���tw%fx�JD ��0BXb�N����V�I5tka���'ğ��\C�RG��ϡ�G��0�����/�[b��K����	'��\�R�����������D�,q��l�7o<C�3:+�X����2=�`�-��Gu��|��Pvx��t��(���x�]������⧟¾�4�J��|2��Y�o���T�#��/cK�?qy�s{�mA~�i���q�i{�;I�t�ƀGAn���>nE�����仩�o?��xM14�R�*ȽI�K��|V?U:.��O��8��3?k�}9�X�r�ܡ��K�t�?[�h�U>�~�bp�i�Q܇z�rq���n_��:B�G�M� ��=�B�&�b��f��.����QCp�G�Rr����@UC`�䶖�k)�KwJ3&sa�X3�]_z�y/$��7m�R��2�jd�)h���Ae��(~q̐=�w���|����پ� 0���a!��I���O�,t�j��SQsHTO�����E����|#g��1|=��������?UԱF�6,�x��|V��5�oWď�+�N{C�O ��"""��3��G�vI,\zO<�\��~N����+6����_����N�R*Gm&ښTJxtp�0�����������ALej��4��\��N�Vo���鄚�r\��fC�--�~�ao!m�u�m���JK[��� ���q���iJ�,���?�3<`rtr@⣗�C~[ZZJ ��W�V����&�u卦8���!���Z��@~L�[�]�;b�s4���n��ė0b��������NU�_r�8�+1����Q��\�5��X�kUp2���"�m�{b>�V"������p4k�?t��B�P��+դ�Dt�4n��`���(�Л��Q*Ȧ��ײ�A	\��p�@�������W�<���w�4���ͽ֌Pb�G��������S@$����k�垺K�u��[}Ɲ�i�&�u�3?������'����(��
�z~BOAZK�[)�"J��[xL��I���s�,i ������������T�����<U�ҋ��Ї��V����dϐ*r��&4;;�junD����Ld8\�jPB���v�A�+���u"|hA��gE������7Aao1�>Z��!�+>����L�f/)K�=v�!�AJ��O���,�W�p�T����`SV�b�R
�_>l�f�{��'?5M� i�����_�Ik��+�B9:����3�1���<�$8\�������=X�ͯ�����P�-�m�W-�D�6��@�g�<���𖯺c����?G�,��?%���V�"{Ž6̺#rQ��yq����(S�Χpé_bO4g����*OlC"8c��Q���!�j��;��1E��*��\h���[5B����L
�{���e��а�I���˾�*j���(:O�7�,��I*�{*�R �d����͏r��R�nk�e����4����	��QX�=�E{U��7��j��.��'����@/ؙ�K�Լk�"E��Z��
�;�G"w0�}1�0h�:V:!�a���c�_�&����cep�8��՛���2kh�[]___�T�a�Q�N��bl� ���h���i�q�о�m�:1��d��k�����[/2ֿ�`\���+�A��A(�M~�
D��j������
.��O��e�����Ԋ.8w��睇�!Q`�g/���ppe�G6����F[��6������m�6�Q��Pg�:��o==T$s��ML��.g�½!�7�:�	�M+x訾'oUxk�N���I�".�/O'm	ǣ��m��=�
_�]Ѫ�{o1�+H�~�V�Yո�[��z�:8��
���:�-�}[���+M�s�ᣛ��i*G�˓�;��Z�%w�����Y�-3'��~8 ���J��0\��ڞ�E�&� �KNu�8b"�����ٻj����eK�"��yߑ��;4�{�w�?�v�����684�F�q�9�e_v(<&��>�B����IY̛!p5<,��,˳i�=�#��o|{4 ��ZAu�jbw��N��$�����^�����G�T��h{�1	���I�UXt���G3:�Zj�[[���ђQ�cM^_�QTZ���TT�����j룇&-ˎ����{��U�ؕ-;����m�d�7��W��F�.��UA��.��͑�� ��D\ϾƠ�[:5=���  �Α��`e��w� ��C�o?zI�P��M�r�[��D��˦�۳�$��8w���Y���n@_h�rXIԓ�έ;ƃ��w26c�Ėdܤ������Q�+��Ӫ���_�D���-o��>� ���t������&.��``?��-�h�Zb��s-CԀ$�X:\��P'�\����#�|����D��)��zz�SU���j� ��`��t��i_���LF����8�G����߯q�s�;r�^yNP�ӸR� ���q��z�����mm<c��,_�Q����c�F{����y_>(�s�<����l̎'j����TҸ���&#>�a�I���C��^��~����r:S����[ uL��~A`F��		�z��7���U�Ŧg��7K��PP�����f��H�q�j��I@m
{�1���ۍ1���X���&�q�϶�$1��j���L�
������J���Ι��by0B[n��&��>�,�E"�>�4ݙ�6GCwg�tXϲ
�)=xÙ �X�e�Vt�����1�Kךm@��:�xVv.ޛ�#����������D�v�W[6� ?pj�%�v6.��žVdzS^s{�8�𫨷)�ŀ��);����Vt{ښe��e�W��T_1�,�D�Iɳ]ץ<�}�z�����1;��¦�T^u�C���w����J(|_n;���B����F�n�j����đC<�>)���G�u�W&#�2qlT��:
�ꁷ��\ݦu �kB��ҋ���q���mQf'��ٔ�'�5`�/�3��Հ�1����kx>'�����5���;0v¹]|��<�/&U��}�۶��:���]�������0�A�������y]�_���,G�=����D���6�����d�A�55u��B���Ə�+����m>|�pitq��cؚ]���1���GH�y���ε5���<�=E-�;�|���\��yb&��N�����tS��:�ӡa^\ǫy���[�9@�#}7�¶')��:���1��&�\�}z(*&����Q��\ɾ���cd�s&I���\ӯ� ��w�����&1��^y��;Ys��v=ֈ�ҹJH���?������F}��]Ϟ=�c�%a�I��FvvN%x`����ҭ��1p>wSVO��{Uu=�u!�Սj���%������iP���_��bjZls�B��(.G0�.�zU-Yx����{"r����]�Vlv0VN��y4����d^D5V�8�&���hz��tѵ"�c�_��c��
<���\8�4�>��3b������%OU���kmi����.�?�r�d�&���@6V]gy���v��g��F�~��@����l���V"�)4��gt�qoHws�D�i�L{�TM���#:�ڼo�ρ��z	lJ�[_熽h��7SݩҗSE�Ӥ�wf����[��x~���v��9�P^�`}S�jZ�hD�i���JF�E�C^����٤�����h^����*K�q[e^+v��߷E�!V֋���߸?NW��f�G�W�7q��gg\�dK���9��W���v�u�^׆�~�2�^c���OW�M3�lM�m�(�
�P�V64��E|r8􊮘��!��E�΍_K)L���b	�Xn���f����?#U5�Q11�"iR&%r%��>�,�m�nF�ش=sI��y{P�������CR���{ͨߒ�1/���P������8�j�G�k.�� �2;�U8���;nw��z������'��1�aP�P���#����)�kn���$>��(�rk%�r�鋆(�>}��5וL�3wV���;{�/c`�֥����� A-�{�ޛ~���ٕ��	��8���������ɔ� �[�qq�������^�;�m@�K⧭xK	j7`��q�\w�r�q��)Ks�-�Z���a1ٝӜޤf;7i������\�M��ĩ̴�L����q9o���6�m�<i}��_pSS���b���Y��~�'e7=w���^)y�ߜT;��h���
R&�=�/�d���D���߁�%�g#����F�T�������V��k�m2D�%�fQ�_%���m:s]ù��K��)����zzzU[�?GG��#Nwu"�,G�{6�O�{�� T�j9|������y>�ϔO�&�!�o榇�7��E�(5 ��Yvw��@���I��;_58vb�]F^�l\F��2��Y���@��d[�{�'3��i�un���M׎�r(�֬�w2N�^U�=�n0ڦ&3-������1KGҟݹ�.��N��1���/�2c����=b�o�S.�|pa _U�����J���՛͵}��]S�g�|7ȏ��7���1�T�������m��ӯ_n^�����x����5����ޣ<~��7��칺ۿ�>��m��u�����ډ��7�1�d掫g<2`�KI.�U�y�z�T֫����`�?������;���ƪPBS���	.X���5��$��5G�fƭ,����@���0�i��h��T��ȕ�b�j���p{�2ngLy�1G q��	�^�P}�|f���J�:�j��qX������*R�Y�K	��r�[R�<>���"M��a�O\��Q/'/�R�����Kq'e�4>s ]D���-���3119�X�W��37��l�rX\⋀����ܞ�KߩJ�蕭4s&UHz�]AR"�/l�`ط������çR=.c�ymmm����i]c��M��珛�9��wq�=�p�%%�B��8�<��2O�� h��]�`.�<P^��,�ţ�W���H�ұϴ�l=�]�a{��S���sx!���IZ�7(����������#/CKf���K��-�k�~(��8{A�H|]Q>�:�RTCV���Xq�,O]511������̲�������.�Wn�	Q��v��G���h$�\F�h�=ijj�z`�|W]]=U�fz�>6���W�!\ⓣ�OAN���bf||jT79���-�C�d ������]7��Iu+����:�vX�"��>�B�����1�)�h�����|�ΝS@l��Ċ�G���i@�������mQ��Tju#��4x���P4�4�:�K=��0mV���u����M�z��?Hdk���l-�,��eKe1K��ҁ߫l�Z���� UD<�&lߍ`L��,u -Ҍq�Q����	�TaS��ȫJ��=�?�_�,��f�����a�dWkv�ڎ�A���ч t'n�9ȜR^i>z��(�Y!uԀ�n�$�`mr�J��gl����I�X��f �}��H¤|�p�����^\��g�K���!��k�/�\��L���Xb�_2 ���]ȨϽ�̴9���@}�w��M.133�;!6XX��C��Dk5L�!�ԯ3H.G.��l[2�/�2p5��D��U�VەURV.�,B���1����'O�e_����L���Z7ZG8��p[饐�����Z���t�lF���O/W��0S��v|!.S�1���E�!L�d��Ɏ�<Wh��kk�����w`;'���K�Ye`�?��D&f�e�	.��Q��@w�/1���,OE�W�JW�!�-g'O�<U?����;]f�K"��CH�uׅ��h}�=i��l����V��.�x�[8��۽��e�.�D������%��� ����}Z�-���2�4�B����|��j�`�Օߕ��g���>|h83�Q�2����ٰ��v���꧹��jr=��J0��R�l�������/--=���6y�|�JfVV����r����W�x��Ek!�����?EN>�ʞY�fe������}�V��d��7]�tؤ�G�N�ɠ�N�?���2�nI��ޣ>S�dd|=�pu�z�����5���}���O�uu�jjj:���,��vU��E�$����'������#�$�������x{jû|��o���f+�p��:���,5�����s�MA,"��w��_�}w�����d	�S��}�w.�=���l�H�Z&"�����d�~���}������%�:y�B���~0�y��(tL\�qZ^Y�x8"�E�!�~��,�(Y�o�cn:	u՗��Td�nmI,���57�����9{x���Q������EB����˟�����(8[�[��A�豱��|�)�� V�����AEN���,?���O ����=�8�&�4�ɞ~�:8���qΊ��cà��i��[���,xg.��x)n�����%�}ڵֵ<u�r�;�WJ��`��l�Z*��"�$�����3S�΂�#�F����̬ �־~\�JKf�k�w�����p��p=?Ԅ�#���O�Q�M)��h���#��"�=׈~�N�|������V��d�lg����*���ٿ�f�_�;�Lm���v���A<	�����uz(�M�W��$�T��o�o����#�55q{p�Ş�k���ZG�@%����!��,w� �
��� ��a]����H����)���T^{,2���������m6.����l���#�SZ�M��0?;������۽8�=i	��"ps;���g;:R�����!԰( �W緁�1��oTH����Q?�|V[�x�ؾ�C�;���CEM�GA���3G�>���CD���ڹ��ǚ��1�"�����U$���we0�+!�ّ��HnTG����O�\�u����]��;�����Ilf/���@T���_rAt*�d�X7u�8�P�1{�r"���҃|�+k��l��\���EMd1��C���������ײ�rt<:�TwZ��B΄�Uq�IڠL窈��(�t)�:/Z�j�pJ9��j��ׂ�¬������K��b5��VxE'#r����84�5���]�L��Q���4Il�p9󅊓Y��T9��w�����t�)�#m��;�;<&�L%|xH�����Cv&)I�mv�gjXa7]��1=��#�l�±o7� �sX��&M���C�ޑx��c��WY��5�ޏR�7m%id��
�!�_kVA�4׉��,��]�u�R�@{�I���x����8,lI~9z��^]qp�$�ͣ���78o�����d����g��Pj�
�K�D�}pg� ��X�"�lr�"_Ѣm�韴T#d��KA/fI�.�|6&Ue�r��%.�T�Ti s�C!���w��t�>�x� ^f��
XK����.'��ܢN��Ng����%��r��n��G����O�U�u��Ύ���e��|�JUg���gz�:����l@����ظx4�:�u��%yB�!.�R��J��T���
�%p�w���e  �i��(Պ�CS$������U�Wu(jn�oܨB�5����Г#�	+�k�������P��wo�(��)��d�jW�x�?�[�6���=cZ
!���F8}��H�=���TO�'$2�z���*����?�VA��@h�C���c@�{oRܝL�۲[�<L��[�譊��E �VL��Up͡� ���d�RS��*#�>@�o"8�t_��1���_�wxr{�@���GY-E�N`j9����N�|��_����Bk���A$t|�j���v���W"�2N��sﭏ��{l��|Drܛ7oznL6�~��:p݌�����A���^J=�;w����+*&�z��f܇���i�����QI�r=(�3�#}Mxؕ���$eh��(����fQ�,��%�ث.�Ш�,��=~�AW���B!�{Y��)k6_<Α��[�ML<�oʿ��ɓ<����	c��>k��m"�KLL�M9H�1��r��P��/X��?2��mq��_�/T0���������WS��i�Ke)_T�X�� o{�.�"�>�Uz�T�U��x��i������#|�N�<���w��{w���8���e�b��pA�.3[���h�����j�k�F14F	 �4;+�<�ya�cV|�%�$N�!Hq�լ>r1��#G�J@ȵﮡ�w��l"B%��^��W*��P�z1Dqt�>F�[����/pT�_���n]B^ N��1!�T	�1R5bbD~-�ލ��j���Ji�Ԟ���C��KX7��"��<�[$���XZ����z�����ݽ�x���vu}*����h,�u����+b���aϸH�i��A;�|R@AO����z��|��O.�ǀ���
��N���N*8�/�����ܔ��}�/�؏�y�n�E.[v�M:,�&���`k�m�k��K���T8�'W����62q�Բ���tB��]���^��>��I�(HT{i�aib����Kc'�Ͻ����j��c��i�<��A���ҷ���ڌ�_�``�_+̻�d.^�1n;� �m��q����TC�,�k&,"��u�������ǒ�`j�5L���[�$ p�^�,Q��
�b�{�F7:ÄVG�_�ɴe0����x���d.��]W�f�#�2��;���,�$.'����@g;�q-��cء��2yڕ���#KgR7�����&�)�%u/���(S�{Lv����l.��y"��T�o���8�x���MpPA29Q��M��>K�����'��u���O	�K@��
}�;~V.�*@>���G����u�'bY��zC��.϶"�(��+M���B{"w^��V�A���KR��)\�ŉ�w�s>��+�.�n|�nBE��'5ϸ�D���8d��a(��IC�|5@��:G���C��.�O䟬�	=1b�Z�0��' �B��s�wԧ�{�����"#����%���qe�q d_4���g��m ���׏��޲R	�)C1�1_��f���r:;;z����U��%>?��zL�bD��h���bMLLd[���3��;�P{���8��<}�����R� \��`���c2�:��?�4�"ʽ�Bt������u_�3���w��ܛ����xo�*��m�WI`�����ﾸ����W?��X�Y(Y���e@/��yo��S�����vޤ�� ���8�q2��-��=����t篡;ھ.G2��u�o�'�>qr.����k�	ۚ�e�ݵK�s�6yް����%�� }E��ؚ�se)Q��~Y��<ʟ/��/o����5^C?�����E��~sc\�=�dt���5��}-p[������(���]�d��A��<,���W}��xh��q�4��]�aF�y�<�|�"�́!�c?����1	�ac���MGfq$�7
D���-�,�W���jk_!Z�a��p��}�˓=;d��W3N�����9����v{Y!3ߢȸp(�:<��\�|�ߺ�"i�&?�zo����z�i3�WXޤ��U�:��-gj27	�s��
5N���ͺuX���ҲM��r-��
BRv��Vʉl,�6��&�����>�У+��̼?ނ&�`#>�؟���||���x�ΐK�U�6��ߨ���T��U�y�m����郘E�&b��3�����qi�e�������_�s�c�>5���>�x�G�i���|AҒ*ш�}�M���ܣ��YA�*�9z�h$��
6�QO��P�s�=xF;�)�ؽ��D�5�{��������P�ˠk��P�;RO��b��=��[���Y|@*+��?�AG��ׇ� '26b��S�znF������A��:MC�ȗ��2'���9���J�繋��1�.aKo�^;Gڋ���șF71ӑ&���'$���W���|�����h�7�coM(�p�[��H��W	=���i�g}�C��D�O�������v�'e���s�jTLw�ܴ�<+�G�E�1,�A^�=O�߂�^"�MV�?�7�&��.Ad \���/�$��Q�eD�s��&s�#8;�0!�V嗫b�e��p��Sz�ެ���)��L�ʋ���wz�=�T������U1�6w{y�]Z���d�n��D��g�r0{����?k�q��ۄW��Y~ N����О�Xu�n��i��	oIy��r�.����/�^<=~��+A�J�_�	�����{�G0�'����۴j\��3��6O�$����& ��Z�7p�,����1��2���9�Jq�7*[���� uѷ	s�R�|D����M�1O~t� ��<� M/�w�+�&=�!�ܽ�|5�7��J�a~�������\���<�p����m�,������fy�ٗ��$k�h���D�[����4��������$C<�UO����m@�u���u}t�<�e�����"�Z	7~xm/0S��c�@��&܍�B�<���%�.�p�?����"�A7�9��m�:ٹl����C���te�4hkA�����2�jw�����)�f�����ku����&�l0� d{�����se�wy(�����m6�v.��.��l3��v<FkN4==�>���� ��9셍���b��h�n��/���q--�|�r�D�â��z�D�q5�0c�d��/�<�K�*���ᴩ4�8�"���@XcA�<p�3C���0��3iqx�IsE�g�A�#�ר���(�i���S��������g���I�1��m��A�_�`�klJ�㦌K�l��70�Y�h1�X2���^ƬX]��=�5d$3j�0c���hӿ��ၽ=�"�C��C�h�h�	Ԭ:���嘣KKKe���g�O#l�.�����SR0 0��g�Я�l��LRg��(yˮcH����,F��i���Z�q��;d�b����<����n���s�ܡ&PP�8�F=��k��o��p2{��]�E]��	�����G7 (1��{i6���_:X�'��䙥�u/�#x`��z�߇o��W������~�;�Rjz|�ֲJR���((-YS�e� b�]�*��/�Ik�n��j8����^���14:Q룜�� ���Ǫ�N���������b,]�1,��#����yӊ5�}_���U���3�K��?S�j	���Ls:"�y�0 nk�E��܂��X�T� o���P�7��p�a�T�SN��N��=�>�Vf4|4a�����L���&��J�86��%�8�)�I���-���y���<��֤�i�0�Y��@��^����u���2��8�<��x��)�rD���e��.�`t���\�$ڏ��T[8�^������7�V3첽������ruNZ:����CM���[�[���cEi&h�"�wê����R�@��uh1�a���7��\p��묢�;&<����G[�W���9ý�u�����d|!]��i꺹r��YGiN��^.�������[,���|<�ɵ���e)��V>��u�v��_��W�GQ�3E���r�
���d9����m�N��n�z����z48v!�}Te�pB���D��=�z2{'P�*R0����B�.JݺAUa�3?�V��
������DP�[��^g��X:�ΰĢ�Mzu�/��ͳ�G߅Xb�V-�UC8Ƥ�#eoOSqkR�1˻��X�?������5���<4�l���v�4��b�'� tvnn��RȜ*�7;܇Q]��~� �b����䛰5;�
�����x~��l$t�T���$��5��坖uI���@'Q:����l�ʴv�_�ت�.0�f�j�@^�o�m�.$<}��%��y�Ȩi�T&!���-�J@սT�D���I
�FL�T7+��'�-ɽoU��F�樨G$ O))�=��~/$Z1hM`������D��P�����2����4���;p�[��{�g����A>1�=i��ۉ7�iFL9�C!���̞Yj�P�5e��L�F�������-���Pn�Nx�GL0���}��5L+mn����x|íb��;K�D2�Ġ�p������F_�Ah��'w_�����Z�T;�������,�8X�,�>p�iY���7n�i�/7??@�t�a*!�P!5�p�׼Bs��?��s�jNf�ϕ�� ��Ƈ�9��X�� L0�J�6�F�����rmu׉g~��"�7R(���nhDۑ/g���dH�@�)#H�;���k݉��_U(����n��'M]��a����]^��'_��R�M��#������]t}��aC�hzz c?
�_�wXH^�.�ዂ_�9��D.l�J@>�/�}ت�V�4L�U�=j3$��&T��,t�ѹ�o���[9֝.��/w�U;�v��s�b=8[�♜7��Q?V	��W�U�Y�ZP�x|��������������?��q�����>��Nc9q����sݜj����IU󳊆�D��	�]eQ6�,x��6fLc�j4�/i |>ln���D�aؒ�l�����J��1a�Tˀ�����Y�*Θ�ʾ��m�^Jhh���H�詈�d�j��O�����R��K��g"h���s;�i0}��u���>z�W�*�H�Ɲ'����h�s�o?����^��@*�%�E�{_��mddem}�&�o���4���YW_*�<iP�v�+���o�"Eg�)E���M����KY�=��?��R&�4"}d{�����7��V��c���(��K�������l2���d'g\* ���)mU�Z ~�����VA����;�Ʌ;3#��
�s��&�����\t� �q��Ș-PX�|���ѝ"��ՙ5�ض��ԟ��%N�뜞|� �u�x���D�d�����Go������	�������{�����5*bz8�eb���R"�0ziQu�����0�Q��b��H�͓�������.��k]u��ǝu�KW���]f~����Έa��tI�fq�'��/+����&����q�44�׳z' ��mUf����0W���!�z[
�H̙��.w��d\���#�>���JJO��xlO���Z\��cߞL𤐽{����W����f���(^ߚ�<��vH-/+���$��n���[�la{�o��{���%r�OY�?�v|�F�?I{�B�;~ ���[ѭ�q��&�4�o��YjF���g��S�r���Z�$��P�2�Շ8Xji��1IvĿ��67Q�t��ͻ6���͓D����V��ǭ;��E4�S.ww�i��?,�Xv�V�*0em���uu�'��}��*� E��!Y�N$X�#+:�=�F0D�K@r�I�Qr�#���pw|K@�Ge�����x�����(!��E�M�3D*#YWF��q�k${��ɾ�.�ȺHH��^��6���5��V����xxؗ�=�s��u��uYm��A�|jt����D~��ƛ����ƃ�\~�'�|JP5��6s�����7��Z�/ �d��]8���9!H����i�'����)ke���	N��y�_r�&�6�֭�mD��zд���=P���\�ᾱ���ǈ�P�ڥ'a��ͭ�`D�_�4#7g<�i��?`-��}a5��>�YO@7����<\���3lMm��`��S���*��IZ�6��8����W��ԉ�l?�	�^g�Ҫ�V�����H�ݙ��sÅZ𑉷1�S�
6���}<����O���R9����FJX;��L����bV��ٚ:�/xM�������M�|t"{���gb&S���te�Ѯ�P��������	B��,a%���<��)Hp@���~<���u�����NR$g���n :��4���bT햹�2�+5�'��~/�d��~��E��
ka�Z">�[����3z)��:ŪkgG�Q�-<�J^]ݽ0*��,��w�����q?b������}ݣ�[�nǾ݆i
j�J��+�%7ا�����Qv0�~~��+Z$j�p,����H�}�zs ���p��f�K����޽E���cF�{"���?�>�\�?C��5�X'�%Fl*���7>|�A�*��ھ�G���������O����Y�:N�i��;o�4�F;@IJ��򒪊	��s�
��	��z����y������״�e��h���f��FFc�N_���fV�~l�me'<���Q�qs�JE�༎x�[ )�1,����ZgbW;U^�1V�Q��H��8�S%�i*|�'�����eC�G�P�p�5�?��Tz��-:6L�UT�;	S�;�۱��)���=�D@�ږ�`���n�-����ȁ-8�:�܋u���~U{s�k�����NA����V'\�U�w�uL%�yLF+ϋg!"q���7�Ŀ�0E��U��uߴ�}��염���vOZ\@o���~�ư6����r9�HzT���k��9����D�I�N�34��-���8��N��NDT���HT9@��&�+ۋ�̧|���Z�H`ܓ�#���-���x
-�b��D�I`�6��{�B	�K����I�3�����^`)-8t����6(�E%�29y�OD������U5�~*RI�RG�	�w�6�$=�&2x�pKp�ޙ�24r8eLz��5�U3Myp�x���x�g�������F�B`�Sr��Iu=�fE�ӗ�I�'�����>���� ��9IK�g��y��6̜b<ot14xϘ��C�[ �Jbr[j`���S9�ן8\�aY�Nֿ�;j���[ ��=�\,�>kx'QtZ������|�;�u�
�R;~�Xo�[����K�"p��b8KMH<���)�K�����|����%���+�Gx.�&�����������zߑ�D�n��`0;���{э�?���F�TLY�_׈�v���>`y�W�������N��:3��/D�7U�_�n[b��zj�RA�g�F�����~���]�)�ϵ��*	l�da~an��7�hTy��^�g6����2xn˸
'im�����a'i���3g�e���`��͖U����$�((ɠ�r��S���U	.ٯA�b�6g����/8�9|���ǫ��n�%�7��9s;�u����V5cj�~��$��R�3B�V8���{�éhu������c�掤O�=��~��o]&�p�'�:H�{�ǡCM�IF?�0u�>]�����47�mG[ݎ��^k�>�UJ�������+ˋ�mǢ��z��q����oC�����v���jfEܽ�+�=���|�у��^��_#z��ܚl�Q��Ͽ���x
9^��� �^����V��gNI	w��ಌ�3�NDssW������2(k��� �i}���_�sC0r���y��� �d��~�5*���1i~�+u0������ s�ݴ=1��u]�z_�OD�s�Q0�y��n����ln��e܊�t���zI�#�~�$�k�g>�� t��ڂ�P9�J~�́Ć�h�2��lFcS������&��c[��.�G�Y��z⹀�Ŏ;�k ���o.�� �l�-�(��d�Q�y�ȕ���7Y�1;�:+&���k�"�V���z{�T�hJ��,{Ȓ�F��1i�,I��Z�~����0tmn��H�T�QϠ�2������e^�m}��V�B3�#�r�1$i�ۡ�=C,!Α���ځ��p���7���ƛT�S0�XS�����*} "���f1j����=@zA��p�P�������:�ܼ6����}VW�ɲR�S�u8r�7/f
���M�	Y�Z�B�ùT۸�C�~�%�Uܙ
���ݾV�v*�l\��G���?U_n����pV�]�LW��y�p�6�y�3��TGֳغ�������}V'�b�=������ ے^��vV���q���F�9\=]��Ǜ���:��*�m!턶u�m`\x�^�s�J��k
}Ѵ�Vɹ����>Ҹe>fW�t/��6`��^U77+�z�DMMmKH� Q���)�n��2m/_;�?��Ư�hٴ�zr���f���嚪��6fe�c	������c9}�O���d������	��P�1�B�U��Л9�Vg�����*  ��K�k�����BTTT_p�'�+�R���+~���+�>�Z���~�*..�/۱��m��-,�L�"��z
�D�5ɪ�h5 _q�+//?�����N�ş��̍gc,�认��CwQrq�q��Q���)�t[��)nf����f2���3^��m��UNp*|�^?��qb�CÛ5g��.���i�c��"~ Bt\��B�I�Ґ��V�_��u�֚j���Ό6�)�W��Ln%j�/%DEC�v��n�͐F���$�.����}sf\b����
3�9�[R���5A����$���GMVI�N���-+�B
�S8y'NNI��z�
<�p�����-���?�N��S9�v��uf�D�;lλ�o5�7�R=~5��
?gH-�8BM�qs�Ip�-����v��Ru�Q���cdB�A os��5]��ocI^7�Zgٞ��V�=��S��:����˛�Ξ�}��+����2$�#�gK�m�~��U��2�J��GU�0��:�����J]����M�2�<��؄�G)���Š��3ζ���BWשX���l�m�=�2=$�K��������@?�V?�m��~Rv�{'B'm�9؜i�!sn�@0U8p�dacc#�B�É*�����l̧	�}����������ߗX6�
�^�����1�R����#�W�9���`��Q��>�=#*��X�c>�x�����b+��E�+�<�:�<0���@;�ug�*��싞�����l�:\[��h�8�d��v�K7t�<\�A>��i6d��q��$]Ӻ�s������J*ԋ���ܹ��d�=]���.�jv,��%]sY����C������q��B�l	���sQ�K�9ʹ%.<u��������Qr��4)B�v��=���n+{��&��2��7m�L�m�3b�ʶń"�E������Sљ��AZZ����z�ӊ����DYTLlع��׌��羅������!c�Y��������jDsHp�:a|����8�������RX��y��́�'Y��Y#'�"?��͔��4�*��x��6݆�I���RYYy���8�tB�����M��v5rI�4��yi��7�_f,y_�/<}Qy�
շ��j�`�׈�/�{��s��9R&{�g]��t)�W&�ʎ
U<@tF�Z�o�4e�!�����nK ��e*_���8�(#���*N<_5S�����g��|����X����G���r��*!^n~O��/�iw���T�'���2�e�pu�fU8��7c�Z��S���=�O��!	��E�S~e �j�͎�OZ�w*���vǣY�=�Y��	Wם��f����IZ�1K�A۪���;�n���Dz���e��ñ[��c����Ӻ� ֺ���S���ӷs�(�3���*߾�da�]�m|�,U����CzfNM�hN���=$�8�{��rȵ��u?�s�z�����B�rӕ��H{�y�VPљ�洵�32�!FGS[  ��H9Q����	ݙ�i����g9��������@v�l�����J�v{�\f��k�.����,,���ݲK��6��8OЁJR�*����2���b;+ߥ���u���=G�Éҕ��m�����RY	��fj��G�~n�z�:��DY	�@g�T�b������[	㑟�nm�\�8|��ƙ��On�Vf��x�d�c�v�oL�b�J�S� )=n�R<e����.η����1�k�34:��m�;���S�vf������#+���e&)�E���ǲΩ[���0�z4���	|��^�_/=i^1�Xvd��c{=����|���l����腶S���ں�Ku�����N��>uW N]%c���7�6��/IS,�.'-��Â'�� �k��1pI�6UG����vO	
���J}�5��_w꽿�� �6/��;e�5�8��ƿ�K2��"��XU��e]8�:Q�xM��'����jZ�jh��j�&D��K���S���G�SAx+� �kڔ�����c8��õ� ��yk\+�[�(�3����N/g�7����%ܖ%c�Wm'�w)�%�g�Bv0����P)W2�nc��Ґ�]wrDFޓD��҃R�h,�C��g���:��O������i��B�,g�be�ј�ũ��6.3T���׉ �M�%�_����<��+��qJ��zR���y�'?�G���E9~��բ��U�cK����������Z)�=I�p*�EX��P�cojaV��M�*�#cD��&"2퍹?M��Vt�aʭ���4�o=����Խ<��C��&s�Ȣ�5�����j�p*����/�b����g�#Rq։���$o�����6���Z $O�S��:�hy_%%�� �~�B	���XP����Tu�v��V<����LIu�]�e�{k�����;��Z�	������1��R��|x���3_I�1���[j^����6����8�*���-���_�2t��[��z���o�@8g�ž��C�8�RܪSe��RK�r��M�S\���qK4��������MJ=�T�+v|�Mj=�b��~#����� ���Wn��hH�H�ib�B0�G>�ͩ�,1v�����b/���߹������J��/$��S��Ho#�7���ܵ��_(�e1P�c_z���+CZ�m�(SO!�lz�rЮ���d ����<����_�`J���N�0/O/}�T�Dv�h4�;z�>�a�"�\/H����jk�}I�w��Χ) ��v��{�6��4�Ѿ��Ѷ-&U�٭-q��tBv&\��b��Bi=�P��5x�[�F�	Ug�<o|z�b&�9��C�Y��G�q�n�|� 7���6]�El�סw�c�r�ǯ -�L��9q�;Y��۝�;<�}���6���Tn��f�M�)E��1�7
��tk6���:�Qɷ ���^�w�#�*����Wk��qK� C��9L�I�=齾��W��s��(~��ĩ���>�zrL�[V �e�㥒t�	N�gcN k���R�#��Eס\L�R���A�����fkv��\%��3>�8�KwbA�Q{���}���_n~~1�cRP�A$�.��Ս�RbЉ�:&�e�\�\�o�x�X��>���K�JH�!�}��Dj��+��������+�6ޝ�{g�s5&N��s�0cf(���hI��0�v�P��]!����I��U��N�vtU+*��P�R}�W9~7 ���XΤ9Tp=!���*Z�/���:����E��U��k3q������6^=�'Rʥ����iQ��<��f�V[�WZ�N���y<��p�:�u5��s��,wy!�f�Yb(H�!o��"͐]��r.q(W�M���5u��D�;�����ۻ���r.�n:Av/�ĺ�,Y�*-����I?9����m�J/�Gu��+VRm���=Hs�R����S���t�u��U�?��^�af��J�c{��:��8	TC{��C��u���#q�Y�'���g����E�~��_�SsM���C�iB�v��2�$�c	�����V�/<���`f��[��E�l�^�����d��H1�Q��aN��-F�X�hoE:�\�Zw��wc���6���'��ϧsm碃<��'�o�GM>J�>�#c�;�����c��DRH��/~����T.���%���M�v@�R�.O�Ӓ�`��cn����'M�S��ͧxm?f�F���/
�*�=�-ڂ��z�@ϩ$x�O������k��0_��z�����x8Ŝ���z;��R��� ��/;�@s��F^d�2;��:=���ykn�@.F�r �Sٚ����,mx�C7o���әtz�t9dc�%�3&�����)u��|����.�@����ka�#���^��s+�B�mc}�54�.��/7�r*�9܎�Y@��<	J����[7��pt���Euk�=6�:�%���������R��8OC#FP|���vqc�y�?!O�ڪ�@mԭm;#��*�E`��oOW����Rd\�./;�y>���zE��)�{<	�X�"-��n�"M��5�#�@��R5ᠩ�	�[X�&�3�Q�����H��"�Ӓ�I�j���M��~���%d� ����Y�(������ ��>��;Y@��lY���C���g�s{���Ar��H��c���Q�l4r
� �D$��}�]K�yʺI���m|��o��g�����S�������߁R�.��{�rP�]������~�y�������4�ב ��ڊ�l�4َQ�i��P�q�Mx��T��QJ�淇�zƱ��yV�
*W��'�Ķ�p�xy�mf�So��x[�l��������ކP�6�!�-�þ�P�AIP�� ���~�����!#M�џ�T�d�T�T��|�뎫��8%ů<��/��%�F̪�[��f����禔M�X�>�z5j����׍�v?[�����p��}Mp�U��F	��,S����m�Ej;�-G��n����������pD#����o�� |t��]X�D2޴]ІK�����O�4G΅�S���~�H�����+S�føĠ���:�緅d:�$�|�8���H���p"����3ox���%�<�s���Rc�ܞ�Q֯�boq�*�Og@��UM�F��i� ܪ��[��xe���	oW�W��s��x�EF�P���f�	�G�q� ���a�{��&�kc������=���XF��B�>�i�e��?�$?5�S���ތP՞���v��]dN�_l'�^p��c�=Z��\�+�;�6�'A b[Ĵ�,%��3e��+��&����)��؅Y� l���i�>�*#t�@>`�,�ʏs��s����֖�ɍ7^��١��z�F��~ϧ�M1G�!xY����G�D��RrZ0�p؝��KO�ޟ��h�
�.�*��@,ö1��Դs6;tW<@&,W��deeϑ�O�<���B���3\+���Ԟȁ���PQ�$ơ\�
1����"������������[�w� ��_��m6�:W~pW����� >���$�Q���$÷��ͳ���?�`�b�l�ܥ��3�Nnr�-�pt�옐����>��=
���J(�`�"ں�ܶ��v�^�_d*>����)H)���\�||�>?| ��%W��~t*����B�s��N�.��[$�Nﶟ��F{��B=�60�Q����[h�`n�AR=����@KN��	�o�5	���i�PF����S73���G	h����w�{?�zw�$;��������|^6��~g��O��b�o��NP3.$�>U~�i�ݵ@C_���j�
�,��7��y�pр�6���=�����s.4�N�_�]��2ͷF�I7�x��� ���2�M�vK��L$���u�Y��:`7l2��tMw�@�I��\2��}�+S~��N
���ag��y��r�*���tSs�����| �Z��լ��
$�8Ri����n�Cz�6�]�	��/Qg�+gH�mED ���!�5��Ԛ�LĤ5��
q���EJ���%^��	���m !��#����R.!{t�����5�[����j�@Y��K=c0^v�b_@^�_rmOY2�^��8M���g+kT�r���Dt4s$�6d��ں�T���:g��Rca�t7"��yxxL'_�(;���d>t�؞�!3�$�N����Ǟ�x>;�U��o�u`� ���)�L��ǜ>��D�u�W,X�SK7�Q��^6Z���q�j7�9=�)���� N��kϭ�ў2�@�qժ�I)�PSξd4�<���q<����������F?J��p6�PeM��v.3�D����Et�L�;�D-y��9���wd�)���@�+؟�T�{�|�u���[|+j`�oX�Qc��M�Ҙ!p�=����*ǻ	vN����1��?���G��n�neZ� a=�s�â��ׯ�Q."����&j�խ�VNʒq�t����r{���G���O��BE �[���4��k��T�j���௘O��
�;i�'�g�w)ֶ��k"�z+�}}�v�Tk��=������v(����� ���p���*z��z���K� RaB'�5�N��]�\�yr���S�?��$y&�4��v߂�d�Tn���S	�����c��7p�����7�ꅅ1����C��{xߤY-(S���d���O#��J,I���צ���|mƙ���$�Drܙ��������'r�b���t1s�k}�'���F�񌇋�68��
�������.�J7�xQ8����ܳ�F��1Vy�H�߯;z���w8h�Q&9M6�<�]�F����k,�-\��@�A����fk9� z_u"��a�wW��JH��)7Ag���V?I({�������{c]{�n 4�*�l5zZD������%A����Ĭ����Ҏx[@���$� ~I6_���V���d�������߼�ww�$�}:K��4-Ѐ�{s^K����L5��6gv��\(w||X$�}� � �z�OD��GN�я���j����{�#傋}C$T#
��\��aY���g�d�ͥ�)�1����NOt���4���lڻx��vi1�=��HEx������IԖ��؈��cf�70�Q<\hO9�ٻ�c�+�̳��6��N�Ɩ]��<���f!�1�"��/�aPcDo� �j.����e���D�\U���JD����E�\`yH9�L��KA?�NO��C˳��=�u7����ڻa�'��a���m�vª -_���C�\��p�l��}=��g���f���4K�����X2;&�Ű>��6�;�ձ��r�-���{�dP��v�b��SN����ꗟ���Y~�<��9"�0�\���>\���w��;[����S(��fw�r��Y<�,�PUJ~� dS��5�1��G��~|愞��>���o�io`8E�L��;�'�k~�w�=���D(q��K�6?B�׿�Zn��L֦����H�v�U���~���!��;��MB�����L�Н����_����IX�e��e�EuSk�W5�X�s$zt�J�Cl͊���4�e1�?�*���:�+����,�P�a��Y�؀���F���oT<�[�ne_s\���/�,��K�җ����Ir�i�}���^�����O �i�.(Oz�1!�g��>;�o�(-d�l�c����#�A�Q#�����ZO�*�	A�$R��]��l=��&)Ӄ?�4��2/}J���{� ����a��ۼ����i�%D��@�,�t��V#�(a����F�%Եf�)�l
�ߺ��@%{";���N  ��h����(\�
� X�]�ͯ��a�陰��&�!�2�D��x�k�9�5x�^<p�_�]c}f�<�P?�t��a�M���W���o�9�t>�-s��\ S�sw�~YD�	�g�B����)Zm�b�@�2&�X���)�i��w�P���<7�G��̚�۹����7S�k�ͯI
�@d�B���9V�Ց��q�e���2%1VY���c�M��1ͷǚ�7�v�c�+Y(�27�/�����!tA��o��l��짲����'�ާS�lz���X�g�(�=Q�;Q$%�w�e=�i��C��
3�jF�~��0VZm��.�)����ذ�5�ʮ$��,��V��0��JeX�"�u�!-�cV��M��:�����CgV,��ge>�<��i��ߠ=�BG���&��ty��f�xG����̐����I,X��㪛j������H��'��ǥ�>n (�0c(��f���9r�����7Dܖ]�$<-T�q�.D�rT
��opE�l)�(p���m���OW�޹��5��u�<��b��, �����G'ʏ����	:(��<�#�؅�<�	�:�?z�m�>�H���-{�E���e��t�ڟj6Dt�O�\<%�:�������{��������k˳��c�X�vln[`u�6&�Fb�HAI��Xl�ae��s�;����^�h��o������g
o��x��f���АJ�{�%�_����� �?�`ػ�$�[RI`k2֦M���`���gxO��
Z�ez迋����
)-��c���V� �_�g��rœt����hrU��3�pM��徘�~~�U!2*�Aj���H�7>|Si�|Ǹgc�0HI���!�}���OT���Ӳ�t��k:�t*��S�U��ƫr_į_ˮnr������F����n�r��Y�}/|�υtGM(]�?�[���R��SO<j(%b#,�@t!xR�-���Y��'!�7�	�����e���,'��A>yش���6Gb�&)�����{��7wí��[�-�tm����'��j��mU)��e�U�1߸.�"� K��C�z�[����s�'�l��;���}3�)�v�"��,:���Y-j��7@��k�����z�!| իL�KE����,�;�\ɵ@fD� t���VhS��=��i?}}r���:����Dc���%�'�Ye�s%)|K˵�y�iِ��	)'y`��V(Ab����
�"In6vp��,��eRe)�-�I}��'aJ�߿����?�!Ȳ��mS�'�'����~��ڕ"��)�u���yI��q�*fa#wC;e��w�V^NW�.�ɩ
Q;���
k��I'�W��
W���7��D�1��H�Ԍ-^�^l*�>d�*���{JU�@��ڒ����@0%$�İݣ7���ӭf6�����ί逪pt���8��:�-���՟��,�Kܳ�o�sJ{���x��5��GL��h�W*mF)�P r'>G�<�<b�3���v�(�5Ta8��;D�@��6�u�/$�Ig����|��e8�qh�i��Z�M�R4�ip� u�tak�;��Z�i��a�UwFk�&X�b7���I"�Eg�Dq��?}���C�a$�CfeS���v�ҽ��R��w4���������ml�Z�����[�A}�cɝG0����X���_)d������&�(��/�&I���u���<���^ڢ�{7���ZsA�l�]0%���h�8�s�P��X'�m�^�-����Wў�Ȇ͹�B-��A��1;6g��@��%l�d�׀z�@��fX�x��vl�K���,O"r'j�H�����<�~5��pl��S +ſ����w�V���4[ �fe�Ti�}tC1D9���)G������;�e��E�����l�{���L��Ћ��|��50��X�u��]I��K���b�\���_��
�7z��n��;�j,R�����<&C_OA[�I<��A��"MnC��0_�⤻�و�ޮAZ=��$%�N����19���ؓ	�ՋwW1�����UH�V�I��m��r\X_uI(��?����+)��*�d�壙�$!.zNذ����N=�ǫh�V��ϷR�������k@���!�jG��K* ���u�߾�$AX��K����f��ϔq�B/�p�ёE������WdK������	^`-8:���xl��K����*��ɔ'8�:!�������7�!_�v���v�'=���F���<w-;F�p.Et����[�����L-�%�''���7Ypv/�'VU6&���wR�!�)M�7��Y/��r��Z�V�\�_�~��?��q�?���(s�sn`|�$��6U�JX�z�H"7e�_�б��5�e��Ӛ�D��;	����]s���G���!�a�P�������f߂%�j|6�j�^p��%��R5�S�b����h9�j}����Ȑ����p��(g�Ō���̼�ю�g���E�ƶ���<�&͆���һq`4q�Mf��,yBt�a��+m�ڶ@�cў�i�iX�h�$�v�3G?���<A����e���'�Z�Z����F�ō��g��`f�s?
��]�� |�6��x�]��a�ҟ�����}���z����I=ˬ �չa��Y��D��*t'L�?>�棎���=I���	N_\~ݘ����v4�eSoHqDZ���y�z���PDU���5t{��>H�\*1����z�	�*"_�����L�!�����>��~��eô�pȦn\�֎)������,5�R����}�>��kI��kt�BV�ɫ9���1�;���@gvh@\�=��(��~��I���rOOʿ�����կ���߿��]�6����C��mY����������5�d&�X1ӄ�'����⥵����ݏϤ�[HNu��ѫu�!�����M�*���"�Fv&��������8><�/5�-l�[�m�x��c���!�g=0  (�*<��X�0`�(%�����(��r��w�xq����|�v�<o�J{�;�A:�/�ܧX�����Tf�1�����U-�� ɛ'ɋ4ck��q���������,�L���Uz�u�PVN�k�<���/+:D��ߦc�Ñ��Z��lO�4�`w++(�rzY@@ to��
Ao�<��%����>
إi�3WK�'�O`���I'���5�a�n��̥�I���7�ă���ݝM���i��+����SЩ�9��ϰS1֥�_����3Ks�*,��e��h�Kk�6'88�� �e�`���NVz�=f��������G����<���?u5�	���,,T�;�N���{U�R67�����6��A )�E��ޘ?�J$E�nZ?)C�e��8�&3�U��E
/��Kr��K��S�U�Kz3�Gi��o������&�/E8<=�b��:8O崹q�UW��`�o���}q�'ؙ+3�����M���ރ��߸ͭ��S�S���~��u.��.�R��k��H�)�륚��G��T��lݘn��[��<��l��+�*��3���=ϸ���g�O�GVH�6�9���C���`���?�p��x�rJh�|���S�h�aW~��.X�)4!���7���1�=�7��c�mG+xe�lڍ��伴gnE�K)�[��rV+�#x���T�\��'m��ڜ<ɕ���ѱ��X��Pӭ��Ŕ{9��H-+����5�m�ޖ��/}�Qqϒ9ޚU_���t̃WOZ���$C�g�_����ض�)�X+��(~� ʃ���)P�?r�$��_�$�|b}�-�Q� �nҀ��`[�nҚ5Β*�`sz6��`{w��{�e�|�(� 2Ra�V�^~0�3�xkM"|���g�,jH�`K�#��g�,�%�=���#���_�&>�A��O��RS&�N�1]�h�6]�zٱ��v�{��D�f1��ef���ᚚ��܂f�F8�>�6���cp ^p*��0jedݖɋ�y=~*��:E��'!#R��}�YҾK}�x}9W��,��'�S�q,�������wwvpڪj��.��~~�M+���*�V��J�����X����1�_�Jg��#�P�S�D"NPWBϸ{��&I9'}N�Z�_��DN�����=۹75�E��X�E	�ã��o��M��/	w+���Oz8��X��'nw_�,?T4����@ҳ��%^`��@���-������V�����#eecf}���l�9��t��T����x��	�Ϥty��$77��F�[����Ҷ�2����[�⇗:�~o6N���$.]ힱ�t��&� ��v�񙛝��M�!9���AU��Wh(�~U:`�)w?���A����K(�"����F�+�	;�9ztfV�k� ���֚9"}�	=NRH�����V'�C'���)�����r!��{\�d�t]��g�|Ɖ�,���sU��j|������M�)N�\S�hXKW$���C�(ljk=��u�I7vxl��@���qi�<��%�������2U"
���03�A*��'�r)y��n�yV$g�0��gF�&��)*vmo�4�(N�����D4�i6F�=��|)�ȷ=�̄��]nأ��T��y4�o������o��g������56LY��z�3��'��\>p�"e���������yR����u�H�ǲ�P�1�����`�Y���o�|X��I.�,�5��O����/s��P\0�F(��D��^dqdw�,&D�z�`��C��� �h���q��~m��hO�BS��C���]g����,�45$���jғ&/E��s<}^M|	^�l�RZ�5ڭ�;Bw�$��	�޿�(�X���iNi��,�D��TN�!��8�#p�]�Ǫ�'�J�.t�&��]� 4:ofB<@���rȪ�����ϖ���6��A�Ӭ��0��Y�#q#���K�����x�s���w��~cc���@�+ �N[�vͦ���.u�9�ۘ{Hm��xH���(��v!�I<��!�"ծyRS��
2Ƚ���.@+�䂍@�d_d�P��t��
�M��-���Hq��Sخ�5f��@�Z<ՏWK�+G:k�ع���f�^�%va�J���$��9�Wᣱc��J��
a�p�)��/H�M�΢��|���X�X R�����՞ڗ6���Z`�G`�%���� 﫥D�OF�þ��k�}C�Pg휳}���w�<��� �RϾB~���J�pF�lM�z��w�^���9y7�u�D~g�J$S�EH&;�z�K}�6p�k&UD��Kb[c,t�/�~6�
��3�_�w���<">��0�[}���x���N�E��b/�����$ih��O��>���ϖ�����u�ik�%��߬nm�8�������p��NL�݈ryY��p�	�`-��{��HQ�C���y@Cx@n<���<�	ߗ|�@:/�D>�M+��C7����#����qH��A�3���z�>�����SV�����_��M�|�gr�Y8�iD�f<��p���@�D��ט�\e������썴]UX��|d�-D�p%b"X����k��D�������Rɪ���t�N}�����u�������V�x��u�n]5�|Yp�VF�8�܏'L��F������i�<>>�}-3���<��&��歧kN�Jwױ�2f�GSC�xJ��� �K�
���|M�lT>r���]�>�S�ߊO�J����w\A2c"�`��	�R3R}���f���`��UY���+��("N�W)��?_�*��
VK��֤
�5��[��\R;u��%=�q����ɹ2]Պ�q�F?Deܻ���מ.��ollB���w��G-^>Eʰ�8����H��t��{s$^������v�*���r��F��o�E�6��b;���$sڷ�sD��cߟ�bV�	��~_[�?��;'���ˑ�?��#ۥH��i}�[�`!���g�B	;r�TsF����`/'dff�~�IN�o�C9�ݱ�l��[-W0�WhO9ŕ)��_%�zqmm��t�y�n�R+x���#-8��u�N�V���D>qS8U�˒0�2�ɥѵ��4�/��[�l���NIc��$d�V������im!UUݕ�N��m��7��^H�]8����[U&�k�`�3���I�Pơ�0-���L2�nVœ�b��Α�O#�
(�nƶ*7m�#�O .���8݅�(��ڎ�VJ���U	����`kF�؃;oi bV�ɘ��{��+p�z_���"f��fi��h��\����yQq:�/uU���p���.Q�D���LW��J����,��_��U��E|$*��
���&��v�� l_��݄�FI	���v	��m�gW�8�� 5�q)�B�����bDMG�S���e`��t���ڍA�|3���������G�y�|��\.w��*ɮ~N��w���R}��}��A�W���\^������@��*�η �a8�������m(�\�;�d�nǑ�vaF�R�n�O�Z����h�M&d7C����ɓ��~aa�YY�i��p:.�3�S�D
q���6P��s�K��S���_�E+�Z����`e�/�/����!�yQ5��5�T\�A�撩4*��>%zIY�SUJO�����������%%%�R��t����T�M����"s��O>G�������."�t#]���HJ����K����(JJ	K/�t
H��.%)�t/���������Ν��<�ܹ���m��+ݜ�U*��ӤU�4��>/!d7���,s=������N=����D��s���%C��͏��P�CS��F��$!pw��N芧r���[+��������Y�v����D��[9����\�A�dmmWe����>����|��s��y�'��<�tg�y���N]��;ő'A��#��њ	�� �N�w�(%���(���TJ^S�����m��$ţ�ǔ��U#i���+�<{cs��r� żK� ��@�C����#V��E��i�F_�|���h�vF�}f�m/��L�~���%����<_��ff��g��9oծ������(� ���2���D`�CP	UR�)����kǴ���f�<� .�K���(3$nB#4 ��?9Ҕ �Y�<3^X_YK͓>�"A
��9x��M+ �%'�Ɉ��=k���ѐ��8G�6��q���m(Y�o
�a�� ����62:�M��xՆ�t{hӝ<"~�g�m��%��fXy
q�X�����lz��O�?��!�x)7h+�u*c:6�����SuU�'�#���;R�o���A�G� ��?t��H��6H9��ʳ�Wҭna����<�?��7J(.�կ�o���J :5~��?�Imy�˹q���.*!�Q$�������U�"la�;����a�u����͆RI����}5933��'��X����zza�W��-#M~���60d����2a�ZfO��5��W�?eWQ�dP��~�Ϩ���;9 I���QOn�H�G���w��z3�=���)������u2���'hUm���v;�-ak�����ηtg��aDћ��Br���k)��̵Y+Ƽ��,f���<u�$�'�,g� ��_t�اII#�]�xj���]��ah�t��A�%W�I�,�4 e�rU�Ҳr҅�V{O (Y8x��YrETP�3��2���q-�,|���W�`}ǧOҽܸ^
��D�ԩ�O��)&2�D|�p���?m�����⽹P��ĽO�=�8jc�?�
}��ocE:ٹ���G�ăc��ui;�ރ�#�k���Ԩ>�Շ��d��&�#�v�ф���|S{3�0��_�i����qEk���8�7=�$�ɕ� ��~�lb��q���$���ؘ�bE�B�Gd$2A��t�vw��*B�æWUQ;=��QaeWi�r��f��*�-P�C�v ��ƾ���6+y�=�b�hSr�-��T_q�_��squ����Q/d���A���K:ܮ Gr�N�7���X���]�{����6v�� ���v:���0��+S7�J��1�ʻ>Z��FrK�*z�|��8����_'ߗ5�w�"kt�aMlC��O��d��mxi>L��&B��Њ��?Z��C��=�� v�߻ᡷ-�~y�f�X�:k.^Iى���sI�G]�n���XG)�Zz��'���;NN�aE�'���}@x�D����"9(��(qp� D����4E�|K���bW������|�0.k.�Y~��^B�H��~�<�¨|�(H���ɣ��7�/��Ytէ*s̟�O��xƺ��+=�`33�A�י��|��6w��!�H��d}X%bz�]ߠ)9+aO�&]�
Ĉ��+�%^�����r��gB��&S
?l���S<~���[�^�?�@�d�|TPƜ�����4| ��*�!�s좭&D�U�����e	f�w
ǥ΍h.��4ުCުH�}%�妡R'���^z���.��	�_�I����D�z#���r�E7�W���{�)�\ �����3��R#9Vq���d`��B��|@�d�����AP߿�v?���IU�7Ӣ�h+��������3�Sv�F(w��y�f
��eh�kF�;��{��J�,_ҹ����%� ��&hfN)9������2E紧�*�ԃ��KJ����������HK���E9���O+�:i�wF	,M��$@P�f u�L��Z
;s����7�(�d�Y��y��a+�4�b����_��	P�a��~maى���Uf�=RaQK����U;GY�d����w��uH@ǉ�v�]��CY�T��-��4|�K�x��^1���۵�=�����WM�$��.M'(��I�U�����yyv�@��=�<M/�aPnq}�3�����Ig�}��ϟ�6���ĵ��{����;��J�����	��q,Z���+
3���h��i�ӺP�=��gl�*i��8x8Ƕ �����z&����H���Ŷ��b��TBDz��a�L����Ǚ
���k��x>�\�z.<������F[�,��Ǝ������b�YCw�V���c�������t��jE:�L�y�\U�?*r
x$Ɵz:%1c��:g?��>����=-�'���$tD��E��I�GO�$<��� �����p�2�"�Pܶ�X����p��/��m�_�����{�a2����Ј��?i��,�P���]�^`���ͫkj��-l%YDBL�k�YN����O���Ɏ����:dV�1��'C�#嘉M*�:�xc�Fۘ���04�2�"�M�iRۗ��'�]��|\ҟ�di�7�Ѹ��jt)�O���̢K�A��5�0��qҰ�Sp~k���/�<q���?���"bg���u�P�yWq��s!������o=&;�]`��J UB���^�O 6����Ğ���Eu����}����U��|������L+MM�i������ע�F��̃�[g���ʗ=�ҘWnKz@����s�RvK崽�'=�h�h7�~��������������qE`V���+�O!AS����A��q�".�����_r��<=�c0drSS��\T�F}'�-4�2�n�;�S�$��N7__Q�l�{����>���˦��*��]H����|�z��L�~Dr��X��̚8PB#�ý�s�A���0�|��+D� �L�3A�5���g��5�}aa�k� ����,/N���NY��J��+)V��6�!�;^��7�L�pXe��E�ǲtX��q�t|o�~�jH�V��"S���M�#R�C������v�V_����!�5���i"�$�瑀ω�1~�l��U�~�qC����B��x?%��٤	4�z����+׻/V�W.�S����g��{k�@J��ʠdg���ɐ��J;��pq�����|���m�т>@zk��e.ψrB˳ ��^V��	��� w�5yrR^(���	�����.���q,��������zl�̽�TE*47�|q��N|Ez��y����m)��e�k�X����R�>�91
�i[���ߜHqw0,�֧�|:����ߟ�<���B]���7�jb��S�I��-���R�8�k%O�;�6�=*�$y,IIh�4
� 8�*��K��r:3��(y��(�LF�F�����S����f�`�_�f�6�]���0�(��0(�??���a6�28��b}1��"��c�X�"�Ƣ9�x����V����n1]f��ͅ�Q1���7U��9�?�f]I��!^�E��^���D��e �����\�2^���	�	~@T��.�4��v�3I0Q�7�ka����0n�����9y��������q�ύr�B���+�Y仓�(F>+����zXbzdjj�	��L�*	����!X�G�/# w�K嗦H�����=@������:׿�V��l3T�e&��8J��:M����]}�I�Q�ۚ.Rbv�P�"_a��[z�lk	�i��|�$�%�R�{����[���Ӌ0�N�v�0�Q+�U#��l�*66v�ތ�V��fo��o'�]@���W9�K�R�����T��hN����>͡���U�w:��2�S���2�� =���Gl����R8�Ks�9����a��EQ��'�z��nP�7���]����+���e��~J����~��	+��@X*���b��̌j�#P��[��)rξY��L�˒py{�C����U�i)����5LZ�ꬋ��`^����M�=C�����ќS����2�/p�,�]�8��s>���i�k �2c�@R�oR��#s�����U�E�S�{�o�]�1c���
H�_��+�<��/�v�N#A��a�	��'���Rv��1�A��'�޺���]N�ԙ��U�t]|��� �NL�Tץ����������{�LE�j~��`F��7WL�	:Ó�X$����"[ת�k%)4�P���P9T���@��a4��OV��vi�Lu|;����t �?��պ��*c�d����~��܈���i= ����0A8�{�+ŻK���baqr0SA	�E�>O�?�:����%���o��_��) ��97U�D�T��!�������S.����W!�,,AA-���a��ʡ���-�s�����L�y�~	����5jS
��N�od��kMh�</�I��*Kj�Fk(�=�׫_2s~�|$�'��!�euZ����D@�=���;�� ?v���~Dnf���i9cy[ Y��239r�f�zv/��[�1��݁_�E��e��8
�
��K�7� �ER%q�"��}���Jo�nE�*�n����P���o$[�/�s�붖Fz��5�҂���r%kٔ���^U���h��v�$���{�/8��yl����KD��E&x�0c�بa���T64��W�P����8�L���A�ǫ����O!c6�O8 =���KO�Q�~��VwT��kw�;�m��	�N0c�z�Q>3E�p=@�u�#�f�}[ΰ������I�N���c@�)i%9��rty^�4��K@���V)��cwW��~��+ϻ��~�кO`��i����c�Ba5�O�"�����z绋��N���6B����jT�fNg8�W��[�k�A�W�߃C��8��"���c�l��F7{�X��I(�3�x����]Z���Y�Ã;L��2�@P
�5;�HM<�����x7�;y�9�c)��j�
�X?WQ86t.��\�~�~ �e Iw�P/zIpx�w�D������2������ȼZ3�#�+Dj�-���Q�D���ŭ�`_8�ց�%w_��'�>�`I���""Z��YP�e��췾'�=�ߣ�{�����07�yF�K�9������	E�Ng�Ӻ���^R���B�tk����7���Ӗ?5�7b<6�!���)Х��fu-gV���!�3�1�}�D9��PX�V'C&4@�O�V�D=
�r���a�S�a�X�V�$�ٜ��|�Za&�MJ��잼�~�?��M�\�~V��''i6�ٍ֭��Z�4���D����I�
�K�S0�S�S�%��Yxy�V�"+5�����&�I׻��쾂LjOAb})�y��q��>��C�Ahs_ޤR���}'�u��t�n�����@�7~$_��G��NF%��;�T}3_AW=�6��OW�L����z����R��}[����P��G}��'�޳W�y\s:��I�IO;7��4}'��᳾�7|�W؆�VR�e{1��Jw&�9W@#C���H��G� ����tjJ����c�֔��Ov�p���fn����T�=9����Z��R�`\/��y\�wH}�j?���U�N��%�@�y)���C6����w�T�\#+J�m�ɽ�K
4�������
�N��~�b'�ؿ3��M:� k=�Fퟔ2�[��J8�U`��k��o[]����Qv�z��vmhh��z��_�)Qh�: �����!IlL����߇�o��J��_1L8
��J��ޫL�̣�p�bX�s|a��Tq��AՎ���{��l,���ߧ��zi�W��''�PC���C����
ܭ��x!���o��s׳���?H�7{p;KCތ�RU�iKL�N�yw&!3h�d��%^MC� �?{#�֣L�y��t\����I�ҵ4�>�pQH���H���9�|�N� u�V#��Z�R~pdW�l���E'���������?�����F�=���hV-��I�X{�Ի�67��D�b�cV�\3&�+��~����>�ݙm-��q�]����a�I��x�576R����]~�/����CH��x2�~3 �	
��rv�e��|#U~���,��H��r|�>�@�#������++*,n�TG1��n�77�������
�ٖP\\�u��HK�,����Z'346�K��{P�T�C�N��;/.���3��Z׊���s�-�M�훭��r� �!�rd�0�ef��I\��]pӒ�b �n��#ŒGY���fN3S䍶�|��\�[{���c����
�~=O�������+N>��\,xdu��Z�Q�R��4���~��� �O9H6�+��?['i�3��Q"&Ǥ���z3H�cI	/�����3,�B�E��FH���tI�޶d���,A3S��.�T�/�e���x���UQ�ˉ�ç����ퟥ�9�~O�� �PYWgW������G���K�����o�������nN��}�1���Yh0�z�5�r^"x�9xy)�U:��S�uo!��S���C 姫'N�6N����Y��@uuV:�uR~(������X�����H&Y�_U�����o��"I�S��u�������4>�U�4ޔOv�N����9��1��[__oPs�tJ����m�t5(8�X$�g��9&>9'��K�!d^/��2��05��xX.���s9[������9��z����W�K��qo��c?��=���N8�������`�\ӁM�����rv���]���U�{ɪ���eѩ�0�A���E݌ȣ3�!�s��5o�W��-�P�^�1ˆW��� �wSk��h �h33���,my)�jSUE�cnBf�%aJϺX�����?>[�-6��y�j��q�$%5u���up��"��
d2��u*��1\�,��I��v�X���4�N���J��L��,L\:���t�O��m��-�_����,	;���R��F�u����kà(���iW��v���]����5܂Q�{;54�8\O��fw� \�U���듛��K���e�����_�������egd���p��*���,��I~_��y���ȸx�B�_`���}|0�0�l�F���<t� _�� ߢ��ak���!��n��u���S�g����LO��]W<ovM�H���W���x)gn�U]]m��Է��i�e�\�>�A��F��O��=�h�?Z-8|�}Ju����Vl.���V�C����.w1���5�>�;LF~�)i�_F�sٛ�3=}�r_:Y�Ԇ���who�>0���\Lpq��y��q��{�b	6�7� ]9���q���	*�~���+!�ĻS�j�Rm��ǘ�"��Y�D��r_�+P��X޸�?0_avј 4�0��������wB�>�݋���ܤ�̵����R�w%�픈�봪pH�;P"J����k~�Yq�M�f�h���"�i�JM�V�e$Hօ5Id��#@�]Igu�)@�n$:Z����㐬0ˁ��Q]�̂����U~��-َ�$J떿.VVO��7�1<j0��~�����-��Vr6�!�a�S��i/�~�5c�4f�/al,���"��⽼�	���j:�j�kT3���M�Mr*��<؊}f1��<$�U�~���jໍ��+s��8b��aW�E�V�6�6��u�R�=?2�x��M����C
�Emu�ѧ_���=%��3.ӯl�Y�l��B��4�ÄOH�Ŭ�u��[Qxs�*�XF�����I,<������,7ifO��T1�=N��F\�s�Ie��-,�����^�qz�	��䋪oP`��OSÑ�3�F�����&�dP��](KF�(���m�cg`ȹd8�v|�`:�7������q���^n�D���@rK!��>�8Y�ڥ8���7��q6r���Z��w9�������z~D"�h^ب�uʎ��ˍ�F}�_T���%3W5��>�q�Lv��
��7� �����ͺ�(��،���#QO)�!_��Fo��/ˮpN���z�Y�F��9d�_�����ir5�"�L*�}�!����bɨq�*WV�s���?0�]�N>2� s
�2�S�6�mM]��ߚ�:3s�'��	lD��S&v����Zf�P=���1�ۡ0�+u�ό�����r�;�˙t�ΣA�3#^Ϗ��OF����
����~
�N���I��D���`�?��	&p�H~	���}A���q�[�b��:y�.U�6���'
x���ׅ�~,��2+�h�@����XV�
�����y�% (}wqʁ����,IU�QH&��UDЯ��웤��Mp����(��X���o��(]]wث����⫊��(�R���G��>��a���i
��b�����o��2�Scs3��%>���<FBL�$�}�<6�ۛ)�����_+�$��h�JL�+mD5���w?Cw�lW.�F4mL}Q�?�~�8�>E9�G��6���(	9?cH|>��M�v�@�MAِSKuI��މ���c� A�T6��	���<weSv�/���Փ'�� �^��4��mZ��5#-�h�tP�-��o�ow`����ԄW�ⷢ߮z�W[��tX��$����vǫV��MLlz���n�F���V���R������Jl���h�d���[v�/u��o�i�]zV��K�@�̄	H�~�NX#cEA�ew~ff��kYk_`q��R�/�|�-<,��/P�EAi�Sp/�7uE�50�T9��M/�M5j!��R����bfH�Qc��pH��i(7e�!�� &S��˨hu��:B�qH[�0M�BYO��R��m�ST1�ԯ��HI�޸�ΐ+A'��O��	J\)�����`:���a�H�Ϋ���{�v���1'����s��a�8/nK,�{=/@��`�4f!����c��M�Y�"D�n�<vs�?8�?Ľ��� X�DM3�مE�39ʒA�_�vM���AU)_j�OX� nIE?�*'���������)ۈ�����y�ۍ��Fl��0-)z�cM��?�L����6q~A	K���W$'�A��T�լ;a6�N�s�[tV����xL���4��E�!��Sl<1��gݨ3��k���а��03z�q�D�̅��7��ք8}0�&:\�Y�eF,S:~������x&QrV7�.��zq�����ܬ(�eA>�"��#͐>�T#�i�HB5u#4�,�n�V�u�6�:�����/p���z�t!4#rG_����!�ɂ�~��z-�u��"� ~�a���r�/�Y�؀p�WElU:K��NھbR R�C,M���6`���<ڝ���j4D9�xjM���y��t�8�+!�l�m��5?�[�|�K��:�}����vzJ�����"fØ�F
��ϽI~ҳ)���y��b���3��0{�Y�WލT%�^�~%���m�����3{��H?�½� M�uN�!<Is�#7��JE! �(1�#奓@|�UݏN���k�'!�]�c�_��DQ<��<S[�|���d��Ӆz�j��J�C��$3Q��r�=���}�w_�EQ�}Ѡa��#��ݯ%//I0{�oH�����q
�v�:�?�t�"`����
௼��F�c9O���/���܃v0�h��x� ���j�]y34 �ϥ�α{	\V���SH�;!>#�,�N�|f�`Ԇ���8���^Պ��/�Y h�v��j+_T@��W)�
GuاoiL�?VCRA����G8x5�ix���M5��l���sNz���
~����>WN�-s.*f\vK���Ɠ�u���%%���b`+�o�- ��]HS�`d~��W����T���D��)el�h�gz��׽癛�?4�M:z{f����4�F���	}}�'�06��v�|��ڍ���z�N���F��^��*�a�mt&�S<�V 12��<�S�/�
}`��AF�8�35=@��b��P�H���
��O�dh"9A� ��hz���^�pE�#=P7I�٭�Yn9g��E	M�7�D���?��4��V-\�}�dH���_�=�
��l/A��|1�/����Î�i&P'�/�t�^��]:fw��^~�b:;���k����9�k�/�� �����^0tZ^����� "�#��i{�[��;���]J6J��O�(E�E���L�͏��Z5}���R�
Oo����l��p���i[y���I�c`�;��Q=$ƥN����ԛBPqbCK温�ow�H=@�zn�ޮ֨#�hs��@jx&IB&=�3�a�����}�X�*��ԭ�QRRo��C�t0���~�l%D���!9f�9�Z�3��a��w��2�nÈs?��)sw�:;-�Ћʉ�����y��v-��O����^����Qra��hhX��׳)���=r2��3V9�~��Ǟk�& �u!N���פ����I�MB��Lx�Wg����Y^��m�z|=G����n���(*��x����M 5��k��� _N�
���u���A��!PX��q� [���b�'٣��a��T9s��׍��9no:H��c'Γ�RFْ�l�����}���Ix��,������%a��ӯ�E;�hZ"���r��8ā`�I�tjv�����mI��
㲷>9�^V�]��SoY�.b.��Yj���l��>p0�>󇉀�)2���(��ӻ���^k�鱃Mj���d��� ���2���?�Ӷ�����Vr�{�C���;q�����g�9�;�_#�g�+KR�[�W�?�Y�����6"�$�Bd�Z�*�Ӭ~��@mo
��؄�֊��X���b���_����Y`B<�ă��FW�j����ꄸ1�)��̸kޱ��V��������h�}b�i,�5<O`�t{���ʐ당|�ԉ���)�i�\Y�Y�����]y����{���(�&�S��9���va��ڝ��x��	KKr���2�=�K�>�v���2T'��� 4G���T?�F��)�zq�M���VE��$�e�
F�_e�rUmi>��~o�pѩ2�$���A-�qߔ]Y)`a�/��L��'>��K�E��Ta�O��P��E!�2��'"y!@���L_��'���y(���'}����;9����؟�/;=���͵�e������8�B�`t�R
�wM�Z?[�U�v��W(�����F�W����@i��!��ay�[�����0=W��q�e\J���d�ȸ�a���WAo�q���G{g��R\c[�M^�>��@o�<�I<1^�`�ɺE:��n�����H�+��cE��֌w�ý��-Wq����V���{%3o�_�P+ao�����ݴQ1?r5$vss}~6�I������bo�z�G����q���_șJWJ�3����ย�GDj��BmS���+@�Q9l�KQ/"ԍ�.�ՙU8���b�5D� ^�"��w�1,���[{5��?VkC�n�Ţ�#��O���7������F�C���}U�҂�E1QM̽ny���C�l���O���%]�8�|��JW�ٹp��E�7������=���.^���my��=N��UQ�B�lTߖ��KcR�Xw�p1ԣ�A��.Ja����pzo#��i�&K��`d ���媟l�gGϭz`F��-�vwZ��b�_�'��k���5��'�fsw�2
�`-�w@��e�ט�$� ��͇��ݷ*J�Q4��l/܀�5ݛ�U�>�����z���t�������(��?�u�;"e	��qj���7(vS)�.��ʶ��:u�9�A%5S�P�bQo���ׁ������D`I�EupK�6���2���4�Jg[�l���*�Q�$������Z�ZiB*�r�91�iq7b�u0<�<�f2u�"uڱ�G;c0J�)hv�MGǙ�x(u�k�o�"mo�b{���n�!��L�gV�]��{A����(�~��p�K�}����S'�*B��4l���>G��.Ԇ�˷�k�E�t���m?m���E5?�S�e��S�[��_]	}y}�e_�jPgG�;����ț9�e]�N�3�'XI��@��Z��(U��Z37���SP6�DJ�8�\V��"=�$!D�CNL0.k��cO��툐?X�ϬCsJ�a���/#�E��݄l�l��vq��򉱘-zl;�LŪM�M�6׻��J�ڂ#��7��>�	V�p��-u��.�J O;p��k����ٛfx-�2o`s���n ^��ڹZ�ǯӀ�^eҕc��73����ڷ�J��r��2ɟ�|�J��?˙�Dg%��KWא���f��dG��3w:��*j,��r2i�E����]P�m�L���$�)KP&f���
@F�^��6CR���L�b�u��l�&|ѱ�V�� x{
"9D^��fG"d=�?�"w�a�&�G�%����Z��.]��mp���O^��=��Q �8��<�uN�؀}�2 l�+f#�m�:�ރ����J��3�2?IY��M�
���ne�/e�!˾ŝ�.84@aw� ������PVM����kO��^�/<d�N�5s�9N����e��O4�Dʹ���C�&�[y�D�@�[�(U3d�	)- ���wgb�A"����Л�o%�����>"������C5��]�N��b���ŇL����:(r�����%+j�,����SH-��_q�g����G�����m\�ƒ�H�tV:�5E���CP��X��c}��ƺQ�UyiA��an�ū#��+��R����u]* �{�: ��3cv2����bTء/�&�<�"�/eP#é	��+��UM2 �a�&�5�vb@�p�]�dB��MZ�)P��������2(��8���'E���T!['���f�ɪ'@I�X8`�{���@�t��A���[ǣ���o�9�	���f����X5�9�/f,/����]����f�J��Q|c ~��۰#< 6�pF�ӂۡ�I&r���ȇo�zxx�DL�Ɓ����*n�@�d/� (��5$��q�b��S����̤s�#�䝁�,��u�K��MB���-g����r�M���6�ۓM�p����7�S�hܦ��i�����g�1iN�fH���~�/�����LlaQ��L�.b n��B��i�UZ�0�i�_��~�V$�q��H]������EIxD\VXԣ����OJ���ǃu���dE"|�?wށ��[ZϢoR�����ֳs�i�7t7�	�-o48%�u����n�YH"�k�Gks7�6�~�)�� �jR���/�FP��ԓ�,��I���c��csĩߎ,}lo�yys�4s����4z��\tw��l>��6���+s{����$����A���!��ɱ���ܤ���9��zUX3�q�.�����_���n����o���2��S�Z-�L��,�%w�:+���O��S��BXi�;�����d2�P���t��X�R4��L�Q�/dL*�.[+�د׉k����n���g��&\ ��Z��-f,Mcv*��u9�l,ǩ"a �x���,��o���Lihii�|}�
�T�C��+U��RC�6d[���\GK� ����1+�f,wsiqY�[����	& �+l�
<�"-��9.b[m��[\��^m��lP�5v�$��;��'������U���M�����	-gK�W?U}�7��Z����BSO�Oa~�^���_�%�W
�[/���w
@���A�;l������>����6�y���S2�Ѽ5�Uv���ԓV���bh]7.Э3Ίy�?7�'��c��O��K:L�7;���,���� ( G��bo<����u~Ŀ�;����Ŋq{e�͙Ok~��avO�BK��yuKy���IɎu�s���A��Ϫ�G(��vC�f��#��a��L�^'�\p]	q�yk�����rצ��W=��s$W�jM�Rsӆ/��q�W����_�g���Gm��Ϗ�Zm�r3Œ�O�g������@���E�e� ����C�T5AT�"��@j�;�rx�qY� [�L��P��+00��u޷���-YdksKNj����,Utu_�>q|� 6��;Ώ�B��|yjFo+��*PR��o���82Nca�%���sF_�G:��#����rc,^��v��r���Q`�s�������]Di�����l��YV^A�#�����[�_-k1�@�{3��������(���;�ަ:}G���A���<ۅ*�N���~�D�+P�1@��o!�o�P�S�!��f��ld`R����ϛc�wv��]�5j����=�����E>r��b�&t֏�9i�[�>3_EQ�7_��46��ޫ��I\��F�Uߜe/����A��7���k�V�����S�Q��DkCC+���9�֫���`��������:����	����� ��5�����ǷA'�}�^�|{6��=�8D����d�,�ۣ��.::�����ͧf��c��v|糭�s�Yǝ��2�jtB�l���1Qr@s�]��'��焪�VA�ˤ��*N��A�r����hu�q�­s���EG6fj�꓏=c���n^CP�8��sٔS�����Y�;or?@k���@eOA��e}�'A��o���	���?����A��M���Q���-�2�m1]�n��Q���w�Z|u������͑�H;K��_��{�-8�J���Л��sް��wD)�!��'yo��Zi���
T�}�&����K2��.�܇����p���эq���������a�K�)un=5�Q}Ae�}p(�)ߘ�zĸ�Ɲ���UY�Y��T�5�C������8k��ě,�B	W_����=�����1^�~�U?�(�c{���7�:�L-~TGw��R��u���I����+#��d�T c6wa�e� A!vD���{@3����At�����ʟ����~�ũ�=ٓ!oU�ۛ�>�@�A��^��~���)u���O[N�8>@�6F��҃jbﵲ�������X����'�N>�X�����0�c���,���wCtV9��7��4j�v �_|Y}-tn����n*������v큸����V1a����G>v}�2bZ�G}�?˿����Ϯ�������0�N+�&Ű��҉*t}V���~�O3�Ker�����'@|=��V�矞��kL={O�Gh��%SdT׵�N>�yB	�0�`�v�����m�T��8�DԚm����S�_887���MU����F�o��!q���Zn�aN�e�@w8��[ҿ�����Y����R¨���vBo�%���yW D�!� �eQ*	�gi�Y��9���l��T��I�>O��EA��)��U����^��7�C����#[ǘ�Ҕ��{e��,`��rL�����t���Y�!"+�ɱ�� ���ڹMQL�B�k^�߁����5)T@`��n�8�'�7hZ�&�J��l����Lwd����r�H�{E⢽7���.�&s��K�;��폤A��=M�� r��H���Jhe^:���s}�A���J��e>M�I��E�P�^��gs���O���qv�`ߝ{��8�^5��z�@�D����nM��R�����z9��^�8�;�+��NǶ�)�2 ��5{Sk��9Tv��sӶ�=��[�B������nW�$��;�x��=�#8�Ы}����@�|�v7AVs̮W���C)�}�ؠ�����#���n����4r��$$�இ���?�k�R���A0/4Ͳ4�6E:� 9�p�fS����_z[母�&�;���R>>�ݱ�'�'j���6�E2���,o���H�Ɵ�O~;F\�_8��3|�8���^�`����ǽ����P�K#6'�r�7����a��а����o(���Rvo�w�02���Ĕ�2}7m�2����i�1b�qT�N�EO��{�gS9_���N�BdM~D�c�E��9��O�F���@|8X��>`j��k��jP�����+���a4n i& �4&�rs�z޳��̱\մ��>�ϱw�������wCYC%�����B��5�-�k�n���0T�ԥ��v ��}���I�߽���NR�M�k
�g�����:���t�X� E���^7'�r�L�f���8�{��wH�Y�q�P��mw߸�C��z[�ȿ�x���/%�Ma�CP���m`T���ז��1�O�A��/!������ 2���q����ivM�t~-%���#���i+�T���\ӿ{�a��kx��lnݐ�c�Q��n��q��ފ�_��b�,�L@B�F<8("�x��P��|,��}���ا���������`�M�IY��,��DN�X��4��E��.����*6sA�x�n�w�B��^��t���	�鬡ʲr�l��C^��*����ܜs;���l|@>���W7b�.�,l.����ZB5�p�z3x�ov���V�jZ��\�Z�<���ޖ�`�O�3�f��A���ֆ�f/�9��j��4��hNLv�$},���-����=��ٜ��k�Ǣ���L�tu�b��ih��ʷ��_���.Ao�%�*[�"Pe�+H��rߺ����U}�!�PO����Z�sV=���q���z��T*�L�Hk�%��hV����~g�.�����Y��L}uT����"�H
()R�A7̠��tw�tJw(J=)�� � �5��м3������`��9w�}�>����}�T2j͡Wf�\X����v2����1v:˥��y��F��\��䢒��#Th�)���a��F���:�������RX֪�$I�y����@���jB������YU�0q&��'%n,�&O�[�qm��YE}�:JUdX��*�|[z��k.�uk�0\�����"�x[���5�0tR#��CW�j�ʭ菊�	��t�'!pMdɭS3'}e�L����a�_~�v���O��ߠI�Y_.��z�i��������f�%���V���pw���:���Ҭ��u,Z�F�Ӹ�|��Y��!���60�L=Z{r(��ߒ�/��67��n=�x�V��4��e�+L��^���7�ݭ���A�o�F$�a�e�|�b�����28����m��>�榬�Qgǿ�Ԉ��Y Z�	�/��H�dE���dG��Չf>�Gc}�\	I�k[�?>�0�c^�R�?�0�%��
Mŝ��F���
;���Z�ɚIW	����]���S[UEw���[�:V{=�A|���f��:H���Ϸeav�XM'����|�3;$E��8j5�t���Q$����l���;-,Oz���(��ߏ+�7yR�_��r��(��=l�ϧ�:c�@ZA9���������b������骛���ֹJ���-�iV�e��k��gk�+�%�oht@��h�S������<�u:�n�q�[�u��߮7o�J���&��W�!�Xٙ��e/��
i�l�Lz��F�W7�y�������
�ឥY���	�_�[�*����5R\�p�f,I�b4�S�C��o��29�b�3�*죪�Ϩ��5n��T��P K]鋫�G/�S�]fb��䡿��gs`��ÏF�5Ė�<F�,�E��mN��� ˽� ��:������v`�]�_��� nR����ǿ ;6���?ΤčVٖ����e{�x\05�1gL�x*��Z�w4��c�m#�96D|hG�:fѲ�k8���mp��#j	D����ԛI�ߡ��EQ�ؘ�i�ո��=��Y���9�moI:�6dI*�ȁ�"O������(���'���Uq��7�/��#s�/�Ф�D�`[!g�肘�*�Ǽ�Y&n�,7�y7���Y��uhh�Ͻ��.������U+��=gF]c%5��|����䣦�ԁ�����x$K�[�6���cZ�Wώ�ל�<-)��|�٪a  +8h����`WD��ݿA��C��[��_�&ؒ�cx@�!���C��5b�/�@kX��Q�*��J}�ﵓ]��f�{���noq�U��;24����U�d��H�E<}���R]�]ޡ3��r]�%�4��^v�����X�Y������9���pr!����rB㫈C`@7�828Z%����y�1���]�2��ܙ��ӧ8��h�����	փOl�O��a��0�������I�g{�p���}	��V1���Cmƶ0�`�u��+�ž���]@MP���;�XO�\~���'�X�n�R����l����' i��^^�#�^�a�ZX"���	f# N��}��*!�X]}|t�"�z�*��f�N��1
]8�����FZ��/� ֨��`@t��A��������b|��HxL	n�S�Vd��e�%%%��t)B���en���/�F��=�4��'�f��A�#|Gw�i��(L|�~r֩}���N�5������槑�9�G�7�F���)>g��O��u[@I�k�7-���x��i�q��x����=�D]4mZE�����C�.�=���4L+�a���9
�6�P���W+�k���BEmDM���X�ؕpx�O��J{S+|LÎ��n���t)e����Yx��s�Rٲ��-���u���G�<T��Gއ�/��[�o�լҍ��1�u�o�2j�d��;�]?��t��k�H+�J'�z���B�0k��u�9��{Ew+3�b��3�m��I^O����@/;�ܶgl�!>�H�磔K��I�A^�(7��jQ�!;�&0���i�a�Z
m�nǅ�Zl��o`�Dg�f������p�z�U�"�O�k��%��Yg&[	b��٪a�����}T���ly'=��2�G�.��z�)�ߑ�1:+`|��tf��B؏m���ڣ#l'��&���l���A�,f"f���#�Uq�[�� \n��4�S�ssM>p��~BG�Py���Y�W~���\D���$����aQ�>�:L��(u.~.�N@������Tzr��<㋕�U{ʕ`ԧ�|?0��t~/��.Ռ:� 	��y�k��Z,��Z��w��D�0N��s)�=iB[.�S���J��1�V�sS�j��׊I��ϛ�!�[6��вz@�����&���7������� n[|���F�����6?��cG<_���Z'���6�(�^ǑD<�j�X�-|3
8����G�^\l"���w����_]���5]�Ȣ�!�c��|�$Jq�>%i��5��%7Eǝ15J��:i��$V= B�~���Hi��� l8��Yny&	w�e�΍'c�!�=�^&?B�"�mw�33�����i��s��g���%�2<�Wj�Z`u~���'�+D��-�q�4?��X��)�I���E-��i|�S%��+�r��`qs�P�vk} �J:�n��k�����[[�/��w�)�����9p�M�n��L�����2��WSl=	.~����&�(���>K[#�SO���]�q�<���L1	^rzg�"�țV|�Ӱ��#��'e�ʑ�?�K��u�a�ͤLҦ�8�7�����J���X�t��d0ʢT?�q�_$Ӊ��Kx�bRw��� ���&�N���G��tMW�<�5��U�;P��)F����b�*>&���il�cV2s���L;0��n�d%Qm�r������@�M��η,�4q��B�_~g�^\�	f��x�V���*�p�$���ʎ��Aq������/a�:�x׈gmEƔP���5�| Շs�̈Z$���zM	?�}y짧e�n���n�� ���HB��׹c^�]�*I�h5�.g[�Bwه��gu.��ivT����d<�0-�/�VuU ��C�?^����=?�'����'�[�����M�ͫ+������̒��{�nN�*A&��'������_�<s�l�}�K�M@A��o ���~�J��e�qB����^��=��y��M��ViB֝k�A���4��_���GS7�e円��<�>�>��{� !~1�H�`�_�(P�а9Υ�ٙ�9��t�J����n����B��è�o�TU��cu��Рgs���7]�QP�Q�訿�-���}g�����|�pSw�[W'�k-.�����I�瞦�.��G +�p�A�. �����}�oޛ �K�R�&���y<�����0kk��[/�D�*	-B@��0���>5�du���$�S~��/�*o��/5g�[�G��BhЭ�h�0�YJ?�tȲ����a�� ��U1qz0���D�$w�����<����.�]2Fy���_ZT�t�t�Au�Bg��oMS�q�������y��7���Zx��z�@��������νd�(�̼�pԢ�I�N�@��R���ɹّ���2�z�1w�2F�1z� �����	(M(���t�h=$�J�N�n�nad~�O����%h�����f7�B�ciQ�y}�adEr0��b��1]�؋�����D|�{[��$���*U6�rs��\#M�BA2C�c�o�\V:v�m�ў&IJJ�� zܔv`Z��j���;�y~��:H�S�ȍ8)=�n�5�q8&4�s��Y�?|w�+K�����ϝ*�V
���:�I�ѡa��F��'��%Z�"��,YY $Ȼ�'r�6�(�G��B���)�f�zv_Jό���w;�������F��%�ЗB�.-2���kNCQ��q
�_	'U���UA77O����8>TyOm�*���S֗��jA�P��-0��Z�F����QNH����\�ék��~��D��6��S��~ܳ�H�����0�p�,@��]$!y�O���R^��%�X3Et�X�l��XԞ��^9͞P*.��o����6o���<iR�4����o}�密2���1�B �-o��|үыjHb��A�T����c��]/�Y!��op�4��rE	k�I���\Ć�2S`���D5����$/��'����/�B�{M>����B����g�W$z�l
BD$8�1�:�Z�=��o���l�u�P��f��!9:�q���?_u���B-�mΛ��L|I�ܠo>��( �����4*���&TZ>�K��4�My�Īc��g�ʻ�xJ$~a������C������aBD�`כs��N���B��L2�y{VIT�,����t������eG�	JV#9
*�a�hG=�*��!�j�qs������-�!ۓ�wH�|wO�
5,Zd�6
&0~����ʅ�S
\��9_�?�&X������<w��uKM�6ۃ�=g��7j��ҝ�M$ 4V�4�F�D���[���Q�6t��'���\W�����;j����ѐ��wc�پP�׾O�8��MB#��J��f�j�j5dy�G��9˝f�س[��=��rݝ��HY�E�rt~��5�J���*1?G4_:*����������p���<��,�ou��Y��*\ �4!"vp�W��&��8#�V��(fm��l=%�~�PK��v����K��D�0{����ie�ת�<���eb����f �H��]��7e���g����GB��h����g�-Iƍ��[T�]�x�@[�R[�W����Sǻ�MoZ�&�7.�����N\�b�êUw�c=�rT��H��o��pKM�$!��ɲ�@��L/�ebv������-z�e� դ�!�J=�{qAq	X}4�Z��O���NDp�?���o�:bj~Ȑw�0��9[A<���fY��dY4�Ӕ#�zb��P�ypV�y�#a�̏��J��x��;����?k��I��R?/���ލ�POc��2T��=�&���9�)j<�1;�tj ��N�?���/�X�t?LR�y��7C_c������z�ʹp��L�ʌ�Ț������~�����C3ϺCe\ˁ`sn%u�xL�n�����Dx�fQ�};p��k��K�j������)1u��E[�����;��)��Zx����^�<�ѐ��E�kv+=S�q���d1�=a�ng�28�0�����	���8��>5���a�&�qL�.��7ޟpӵP(��3ӥ?+T<W�B��6)x9u��H�CK���°�u�6ܽ	��z�����+5�����>*[�ʾ��
���%��g1���y��s��%U�����<��Q�V��(�{~6wx��dόώ2��^[&s����C�Ky,��|p�����7?,Rˬ�g<m�gF��������n)�9h%�� q��_nU�66y���� �U�޻��е��93|��]>�A6O1͎�n�9e�Q��ez<އ��OE��3�kAXXT�o�2��9�~�OǸJ��W�{oy�N�KSML�!؉b=}��S���KE���џ��@�gȚR=n@�x�����]��{�{Κ��A,�>�&s��� ��O�7;�}��\����<��,��ȉ����D�j��9�x㣧��i����h\�����u"a��� �(��V��R�������1�.n�� @c�}?c���H����@ �������(�l>B��bPq��lg�툱+�8�����)K�R=�'9��K߅���wZ�B���T����J�>�xy71"��w11̂�7>�~$^_��j�BG4w��3��*RE�|ӈ�
���>�χH��b���^�Ւh��`��M�PQh���@�]ԗ��G�p5�p	�$y�D����sx75�P�(9!s�:P�|N%j;�@��|��,Dx�Ӏl��u~L�?�p�T�3Y���/V
��q����뾝X�Ϋ��exϸY�� �R'aQ�;;�Bl�&���g���6��,�۞�TSB���G�:wE=��i�����,�`ؐ�T,�#ۯ{�8���d����\>���ج�Up�b��>�ي��ؾ�)�38�w~V�GM,Q�=���S�.��um�Xvi_~�;`y�R����x@>�z---�!L����9��:@&W���r������O�i����t��Yg���E�AC���RNyN�.���Z�lY�][��aZE�!V��2$R2fJ���2�%��yC�
J����w]���sEP(	
Ձ�ɻb�J�a�q��zP���-Ň|��� ��;��Ѻ*�"�^���Fk���f� 
d��	�z9s�F(�\\\�"����PBv1(�=i���<�[['���h��X?!�`�a�<�nXn�?�+��gI�ob�ɲ�	Lg�Y6�����k��s�N7���6sc������+�v^n��!��"�������K�����F���	�����H.,$us�'���$��y-�$9��z/���t�u��e�K��,2�GZb�jn�_5���sRF�?X�ϟ����fR�;�*�L8�_Г>�w�\����ͩRx�pM��)��0h���]�<Y�B�N)0e>�� �sq�Cn&���b��9j�k�9���&,ӓŶu���#�?�Z�?)��P�+K�w�j�v����|�Y�Uk���:	��A4�]���2r(g� ���~�1;˩����)z�p�N̅�U4�=|��#�Ȍ�V��9)K.Ki�o�j��bS�����)��-���و��ʉk��lnŮ�[p.���)�T��ц:@���O��]@c��Y����������V�]*��-��8�)�Tio��K\�0���!�������}E��w��=�j"�W]�������?�<�y�(G�S})���9��6�&>Z\������&��J{=be\s����:Gs�X'{�F�^Nϥ���\�V�~=g<��w��}�����]��	F�Z�(Jם��"�c8)��w�Gq�.��۷fmEOWH\��5��<Dx��K���id�i�`v0ȐH~�����?��^k�fu?;�������5��;z�9��b��\����Ms�w��;N����Q���F���Z7�Nm1.�88m��E��ǭ�p� ��z\?N��csmqX��<���pԬG7�.
?��3�3�!/gý��F�)6<�B,����:�:�%���6��4;o~�q{۵|�����='�]e.�����[/B���F�����+�7�W����D��8z~��P�<"F�{r�E�L�^���?��,�"B[V��M���k{�Q|_v>�4�=Y
ן��K_2���G���⠹�����}�$�<�9NgrҜ>�|*[�8ⱗ���\����h��Y󉵰�BK{,�z
���\�����{X7�z�A��9G�-wU�)zF�֪����[���VG��n}�efu�Ё�;(��B��!r׹-���հ�\��s�+:!�,�*V��Z�N%����qxo
�hJ4�����z���L.���8]juGM��ŮL��Le�y;� O'J����~\�-�y҄�*kZ��XsXY�g���=��_dJ��i�E
�������<��6�r����r��T7xQPNFf�Ƕx��k�y|�~\>�{�%�}��9r���}t���V�413�;�Vvo/;��Ȉ|�	vV���Dma�	?�,�-pk��3)**�\�Wr�I�#U܋�{�Y0�GQ�K[[[?�>I�������j�Uk�m|�`��#ח�f ��q��]�ⶦ	��Z����t��_�IJ���#z����J�۶Y���� ���%w	0X[q��ȄSF��ԳW�"��x�'�
v���������{�w�4�x�t���Z+猴ܳF�}cw{r<�V�*3��`�h8����W��ӵh���sW�k�-��M=���Zv�+$�NR����j�rA�	Loc��
�Ə����(�;����D}���3k�Y�
kMp1�NY=llB^Sy�Ū4�en�E)���A��Ҩ�}�	q�kY���E��N]Lk�X�l$s�.<8::��(����=���K�C�������q��tT9M�"�*��1aĈ���G1/.|�cɩ&��kcm�[�X5�F���7p��+��\��t����7:oȟS�?T]n���'
(y����5�d4����ܖ��C�y���g�%��Gh� 6�2,k��۳����)��nذSF��K�x��,��H��\�� �.�l{�	��p���H�R�~n�����rlIRNG1h�7�sb�+��uH{���I��v� �de�`T���j�6n�����Ȥ��7_�܆4oA;Nw9���Wz܄��g�ٚK�Ӽ���y�Bu���e�$G�^4.�"��."b�%B��:������S�ݯIVs̽�iim�Ĝ��bBk�"[��O�1��o1�I�{�����aHwq��s|��-sG@�3�e����cL�����Q��05��u���N��.#P���3:{�����L<*����2zhХ߼N��!�F���\����x]����ɇ�|�A��Lm����cqB�V��bd�є�<$����$m�I���d?'����&���"j���`��1����OQ�K�`��\���%��M����s4���Ǥ���4Vc�ǵ--���r�+�Q�z��d���wA`�Ne@(�7ȑѡ���(۟%u������KZ'����Z~f��R��较B�x�s}�c�s�k�"wj7�J_Ǧ���.��/�kI��STId&|���9��u�J���f��\B�T���v�J�DAþ�yƤ��j� N&�ŝ�^j��NO��p�(w�{���tَ3^RCx!�������U��t� ���q�'�X �2p$���~��ӆhU�R��Ɛ*�O�efZ�t�W����i�4꨼=i��b��@k8�E"?���=<�*o$�N4��n{s��Q�mM���K����v�ræh����d3U��.�J�Y��A �aB�/�;�9t*�c��էMLW_���Z�@��n�95!*r��D]mm�|L:8�h��V�o�������-��~h���$�V�}���͌ڄ������ח!A%Y�1qH��"��rЫ��gl��S��Rp'���8FhI_ɍ����#���H����Y�׋���8�L0&��q��G�B���u�L�D���u(�������5~���7V*N{<���*I����8)J��4�r?ܶ�bL�IEY�W��woV�����]\Ȋf:E{8B���,8&D���݃�7�,��D����o�~����)u[.�)�c�M��4�K��"zB����:H�4YЋ4ϲ`N�����t����ͯݖ~*�z�<b��5�J��ɖ6��-��/RA��,��g��tw��d���o���S�L{e��������]��ZIp�<�&u�r[���Z��y�ڿϘ�
&�~��Q� ���.�۝2B�{�\��� ֖G��%u~��@�lrÞ���XI���×&qbP-��A��������V�(��[ac��p�+�"�ֱ$X�.�+>���)60�r�c����j�V�l{�Ԋ�$ ��<>�q�s#��:� �ͬ=�!����m�8���c�߬��_���?�t�#��j���~a����^��гB��;�i��v��?z�x#�ECM³syL���m%�C^��u��B�?���O>���Ů	W��0��n�E�wH��_f�t��
���.��>C�6���M^9dW�b�L�Ѭl��F���<N�܃�(�El�'bca?��a#	�"^5M�8ڥ�����8_�nv��E���!���7���l3����kK]�q���y Jje!��f�/���=����u�Y��"���#�F(ϲN��g�``�FX�"�A���|��孖��J�v���0�I��B��i���'}x�gX��E���h4ѡ�j�E���4o�O�rz��{�������@���r�3Q�)5Q m�ʊE�W�{3�V��[0Gq��0ԕ�a�R��̓
N����q';R�U�~g쫃C6f�GHG;��(�����Q�~W�.)�p����?_h�O~���E���`�3��ˎ���Q~1x��=~����$HLg#��zܞ��]�F�q������h����tꤨ"���^!2�7M�%1$�Y�Fʔ2š�����z��s��uB�}���6��qf�o�����:IDt��D�x��l��2_"���FV��*�����7�o��z�d�d_���j.�d���I$���"���?��J&�]����ڲ���uXGJ��j}��:&�ydV��6�QuM���Gx��BC�=l��(���-��hS��2���9�yD�̆�6I�͚�4���| ��P�ըOW�D�5��ߕ��OT	���Q�]�GW�悒�N�0�^hŽ���9����^�'!�������B�~oV[n���?g��*><��q~gE��ҥ�1{�WW�T�<�@+��ot�
�|��I2G[��Z���d�Li	G���c�:
'
3';���Z�$�>x�V�;�����| ����\h��lڞ�6D�9����R�����=ȎS77��e�jq2�Of��p��ޯ���;�d���o4}���K���G"�M�3.�{�a����=z�����F��}����8I������j�h�Ar䍻�����KS�Ompk���W��Ï��D6[�%ade���Q_���lZu1��E���]�l�����w��
��a1��؜C{k;�v���J}��Y��_ǡX�ѯw�$�����d�ū��B��g{��J|ۀ0���o�}QϜi3���Jo��a��!N��r�JD�DKR�|����V���Bq�D�Yֳ�jɚ'>����	iY��K�R0X����d��~|R�+��ڿO�%|��s���}ٚ=��y� �?��G�c�i������X�(M�p�e�f.{ؗ��(�ٰt��><_���]1,!0(����� �X��ٓA����?�Ur�=O������Wz5�nz�z.�@��v�5�]!�a	˗4��N�2��)JN��RO]TdO~�>\�A|�so�����4��Mq��,^��]8�>΢�f�����ǂ�$��s�E|�zm'�0�S�]4��g��7��@������l�K�ċt�'�v��ݶrd#��j.J��a�bv7���+��sr8��	u�����ڸ���1���y~@U����\6'ɏ�� ����Cw�s���0��5S�K�(yv�o�ML�}j)����e��+UAn�맫�ǜM�+[F��!;k������6*؟�`�p��B�L��*W��+�&��p�ϯ_�C�*����Tq��ClMt��-e�kϤS��1\T[fwgtu�c�GH�"�J�(:�C7���T��W${$�y���h���A(k�h�rB﮶f�A���矍Q�¨O%�a�1sa���`���c����?�um>��9\��;E��J��*�Ԅ�2� a٦��)R�'
k$v����e/��u��62r�"��P�:�Vs�	�FG$2QQ�Y�i�yr�BU$E:!��Q|f���:]|����s��f�����q���}�u|����,C������}zU�s	�\��9��m/J|*�����j��(6|���e�_�����Q��U�ϸ1O������_��Z�t�M����7��X"+�CR����s7�c,|�t�*�"�^���ǽ��X�K��l{�|8W���i�`��?6�rP6�u�c�6C-�?���7�.��υ!C��vm��	�B9sp�Z�b�q�'��� �����!�+�ytH;|l��*���һ�4)�N�w�ӱR'	����[���(ɛ�����z�K�O��?�@�`�t����'����>U�Sy]8{�ˍ�X@Y�]��ׇTmΰڊ�/�ܝE�y<s�Fv��c�=���)��- ^��9�b�e�� Y;��3�u�?u����|�(1s��<]t��Yg��_�i�O�]KV�,��"��7*d�5�?�o�Z�"C�{Mf�+�US��٧dh:��(ج����XA>����,�7���م�?TeN�I�G;_*!@\QKi,؇-7�l���w��ͦ��q�[H��u�P)��Y� �d�d�� �0�L�=�d�Ȟ��m�8�����r���~b���!!2���=������_�+!�g���oy�92~})����M��<�^F/�b.37������	������9�a����#Ł� m��Ϊ�(�E�8D\�S�U.��*����mۘ��т��N�$u�����ع3�y�P6@���)��om��ϫS�d���Hѕ�8�W��T����u��q�iw�U�QD�u-g������!�໷'&�����$t�g�~�r�l`S��w�f$�p
J3�F�g�녀�H�c�G������v^{���-n����rm`�������t��)s�쬎��xAL&��a�N���0>��̯������p���nVgK�t��%#D���Ƿ^_v����h�����/�J-�s���#�|r��X�{w����.��1��͟�h�W��z���e�d��M૸��]�uc�
�ɔ��Vp��u���֒���ЧJ�eɳ�h�������'���u;�0����Q�V���ΰ��	J�a[w������u��<ʱ�Sq�ʩ��(4"+����wg�DRl����U�`�;e���k�{���x�l�{�I���I'듨q;3_��7����鱒��4�(���j������!{=������%s`��KTug��-�{Rњ(�����p�=�����K�pX���j�qWA������&��Џ��Ct֫�~������h�<�s��9� �H�H.cnV��>.!� � {	7ec,Ó���al@�3'��R܉�;��������E,�b!"��X�ɛ���\-�o�j��Z������=<J���I] y����!YcG����9Ӳ_�ON�a [>V�X�L���+!��=�	�(U�:�p0�;CW�Ҫ��mz����V�n�(�7&����v���{Q����u�D�1�Cs���w��(O�C�c�^A�չ����?��;+7w�\�7oBE���\)�D��2%�s��n�5�A1�l��:
YZxA���c�Ղ<��7���ڊ�w��C�T�5����v^'�d�+l�]%O�sS��ս�P�ި90J����طB�N,�h�vɳ��K��L0�<�~u�>��y_@ό�5��$�����%���+4]�Ⱦ�݃R!��F���Ӿ�\�wD������6�����]�/�����17d�E� u������s����Ƀ���Ҽ�읍rJU�H"����1r+�ą(�8d���m������c$��͖+����D�¾��R�T�2����[�u݆+�LN�H�L��Jr�W�y�+���>&�gVZ}%?�>�z�\Dn`�N�2����!��A#��3���G����\�q�/��v�J�J�p������zȶ���u'�i�������Q��a�������j�z�u��}'�J]��l����[
YZr{m�+�]�h4r3U6ڱw2y�vny���	�Ő��X7֌p�<�����o�!{�r�tn��9X�`5���Qkv&)Y�����XA��: y?�A�o�,�,�3y7��1tE(�U\OM�E�[A�^
n,�����M�K�(>�P�Fz���Z�鋮y͏��5Lǘ�Z�8���T)7Y����O}%����F�60�_�3���V9��skS����g�m�D37f�-qmB��"ĆZ��_���.��"z����%랥Yi�.��^Ail�a����F}��իv���\;1v�e��L��o�!����Q��v��y��d筕�7�z?~y��&<|�{������Mw0��	$����M���Ȯj`_믁��FA�k�����3t�OA���e�(�w�;]y�Ӕ��c��{`692}���D]� J��,	 �DX˹3�f���9��N{f`�䌾>��-�������F�Ǒۻͧ)�{-±Q �����Z;+��rW����o�g�R��Nv���s� ��YK��A��w�*׫�����D?6��S�H��{��{�%d{+;��z9��m�t��U�jd��������-��K2'�����ٚ�p-]�nİ�����.C��㸯�6<�_=3�?O��Z���ע��ڕ*Œ�
=ht��r�-�m�w�p}�p��z-�p�CWeJ�j�B�����d`����ܓ��:qC]ݟ3[�����X�e4�o�oG^_ӓ�� ��s1-xݰӐ:pxprJ�� R�0�F��*%�q{�{�S�����uh}g�Zn��{g�O>6�hiߓ/��~�0\!�96c}i�������*�	�LW���t�?B�z��;q�Ĉ��~݀��\|4%�5���Y:�vԧ��s�Β�E���^��U�[ݐs,���>���v��@aY03@e��4U/�y��j��jb ��r&_�o�~v���|���*`�᪖�}��BV5�ǤK@�+��k�����58' � �9����d��pF8)�_�_'_�Zε��-�A����s�Ng��^b�O��Ԙ��^o__���lM�4\ː���M�D{��5��z��L�Z��^�����n]�O�{�}��`o�L$����5�`�W����E�H�G�?��z	e����|�(�h��	����(>cuG�HoQd?�A�����n�+���\C������������v��n���Y`�۟f���W�ep�'�RÒ�
j��>j�{b���f 
�U���N�Sb���Q<�T���@�k���F�QƧo�/�;��z�Q[P��j�&�>6ӽ	�A+��e]@O.N�h��` 
y����������p�� �ba6����%�ݔ��4��/E�ޚ�
�z��"���5���WjL2�˛ϊ��d5��\Dx��˂��a��1G�B{������T�H��j<��0�8D���4C��@�Ã�/���9�쥯��1����z�����q�%#�m���̜g\��:İʦVQӛ���w�*�%�	�Ś��ry yS�J��xD[J�^���Z����Kv��n���"�[=*�;��Sc�W����k9���~K��^�0k�O��ռ���1'��1�ҟ��Ő�J׬�l��k�ix�=:8�ŏ�_y|��&E�L,����(i]Ŝ�kߖ�䥩�ܶ�6s������;�� ���x�0��/������y��B�l����:�ɆQ=�Ō�f0w���,wm�"�r�)r�ss�KU%����!U�?�����_���zQR�L0�v�s{w�uڻ�%����������]D�jY��5m���Q�/�^�D�����(��>��S��ˠC��:V��]��e0m�,Y24R�#�㔉b��F�����h�G�yO
RD)����1�^��ॕ���k��.ׯm}���H����_�/"bQxm�JMIᗒ�nk�c���446q'L��1Ȓ��FΫ4�`��j1����+�S���Oa�L�M���P�Q���/���0�������R-U.!j���/E2����{�x�5%�`f3S܄��u��L���͛�<t��ggg�|���4V���]�t5T��!�k�A�νϝMv��u_)v��^���~>goP!܁JYu�(�)����[@=7�~�;f�s>��bv$��}��Ȕz�?�^�G|���#lT����X������1!b�U)D��ƛ݆�hE�0$�>�X�4Q\y�x�\���Y������ޜ0sC^(<(��˲~�n�FS��S��G+O�4;�{E�E���Y׃���"R�Y�ec����`��_�K�fu��Z�H�)R=�s�M������#����r��U�]3\sv�秳��z��إ
���-T�-���~��� 5L��[�o��/�����<�I�OGd���(�].xܺy?F��;��m�02�G��-�oaoA�Ӂ���w�ߍ�+#�n�����-"���]M��&|��!ZvhR�
[.^r'���N��Қ�����Qi� �^�������s��Wt}h9�Ӷ6�k�� <�#��3ٸh��������%�}5d LR�q���������r��o}*��W,\��:q�?�vK�$j�3v�9����"Q��_#�|a!��t��9��
�U{��_TT���,��~b�7���ˆ.;3����:h$�B�����tb>ӭv��vfS3��C2�P!�!���XqK��r:��7-Q[�/o9*�"w��ܝ3b'5R�����K�cm�5���9�_��:˄ֈӃu�3��u��~d&�rl|�`�b����Z��mKrwM�d��F,����mί�:�Z��-*�c������=O��ҟl��n5G&���k�O�i0ƕگo�R�����j]�fn��+�D�`��D��O�7��No�j�>�Mi���c��~���P�,{$�$G�Ǌ��lG�
��������Q�&78{�P�q��͝��{_���~���ǽ_���9^����K��k�r�R� 4F@�
�q�c6���e��j���`@�A��/�d Y�㈆�4x
�'_f�����+��ѷ��R���ܑԢr�Z-.���6ǻZ�w^j�+|�bjsg�I�� +"��٠1qgh~Y_$��w��=�lj>:#x�i�3����p�����
a=r����awF�!P�٢��Bi+��x�bd�z#`B�\t�X��U&?:m��djju�"�t�w��Uϭ� B������S�OvF���rNk+/oA,��o�7{�AU��v=F�)٘8>)��Wy�'"���W��eQ���6�堜&0��("����k�'�^=����m��^N�`�5��t.�ez�0}� �:�1�:��vM��q�`l?�z�3&���b
z27;�U�~�"t������wL7�	?c5��h�Ey�5���]�5�ps�q�[C�7�z-88�{@`��N��()��F,qᛰ_p�&�f��t����F?p�)۬�v^��%N�
.*���@=%���<��b[�C��w���(��[Q����ۃ{��8����5�nL}����ks��ppt[�U&�߇"BF�O:vUPg�	����m}
�=xx
��M߹���Y�0�{�]w�����'�@�xi%��^���3�>G��m[�\��6���������xT8cUd5"0)���OS�P��`OvΎ�����ي�56O��|x���9�Q��+bW��.�c�Z}����Ib���N۞��牄�y�U�RW�D���Ү�-�L��ɺ�67&	�
BwM��f�P�K#;�K#^T�.ff橄�׎yE���m붌���L�L�sH��;���Ҫ�G|�K��\���kB�M��j��/� �c%��͡���|�Z|�c�f�G�e)�<��p�������� ���[�%�r ��&��K|�tPI:�j9��}w�7���kH�{������ĕe���8AO��%}��x:�DRR�g��v��K�e��%4v-������(4>z\�#���r�bp���q���?�?2��cʭ;w�K�t���p>:F���ɪ)��4aq��G�D�/"JEg�F�5�`1O��u����2ɼh�\v���9_��
jw�,d\q�U�n��;� ˙)��CL��ΜivKл~����(�2x{,�<c�r�de�c����|��K?�M�f�S�l!����I�����х���_�U��N��~\)N0*e/#�}G���}���]�"Y�u��5�rR\�	l�u�ǡN�j?�5ߛę �`cs��U���xK���3�h���)/B&H��昂&A�NU�	��z�6��)��Y���X���JF��N�_*��Av%??���_1A�ߺkP�X�Y�]�*ZhR=����;�|S��EsƢ�8[���]�hp3�̯��f8S�Z'CW~��X`����fDF�����y��:?�#y�^�L�F�L�ɒ�~B���?�<����m�3Xkc�]6x�}v��' �:L�q�,�M7��^�*±�����)�mb�A��W
ȹ��0�(����Oޗ#��s�J������#Z�`z���A;�<6~�)F�*��ڜ�����$� �v���L/Ek�!e�Ҩ.{��ٷq_�B����	qa)|6�`ft�:iO�}�'%~>���� E����ű3�+���<����WY@��O�>��6.�Oz�7�H_��}��^��{�w[$����ڟ^�Vq�u��_�I�R�DF���kE��CQh|�����QL܃���(c>�B	s���+������ ^����܇Z��~�~4���S{`�E�(�#*t�Q��ʢ���^&�y���d#��El<
�i��xG�/�Z�0&b�_{�����U�1���h;�#&m{J-�Aޟ�,�M£�C��J.Z�1Ny
�8s��$5՞�@ϲ�]˅T������Ś�����(�V�ᜮOw������s`����|�n|~��7�`�8����cR���U����^j0_Z�TRZ��un����H�
���S��҆�k�)xa}H?OZ����f*��67 �ޙ.�B{y��x��r���:Ϗ>p`�!��:o�L��:����*QK�w�h�����[�_-q��U�!�HR�W� ��C�0޽�3���?�xN�4��.�����35�� 32�Ѝ��O�8�)�$NGV�\@�5����U������5�^�k����,��ٷ��~ʘ�5J[/��27&0��ǥ2��ON�+X��g=92B"¾s褂(�>^`�r��*Z���ǚ�|������$�ӨL�K%𶼾B���"�U�.�3�b4��tKw�Z�N�򭩈?������<�v�4���`���qm�Qz�\��z�����w�6kc����z;y���L�-���.��'KL�Ψ�8f��Y��Z�k��*6��������.����;��AmRW�3/58��O���q��$���V��&1q
$iM�W2�R0��V��1
���,>@��Z�s����g�/��E�·�*���=J(g?���#=b���)VJ����ˈ�z�nP��;��zqO�����U�������z����_(��1�٭�_�:O������?��t�3(�PB��.�?�@T�HD�&2c��R䂞R�*|~&�)��*h�\����߽�<�<"6T�����[}6M�E�`g����:`ܱg��9�ò�,�m7��ŔlP����u~7]$��L�<,����3!�BSZ���0r6�5�)�L7H�!:T��������gTA�P���CËY:�_
�Ҏ������x]�����,��)�/���WN~+~�+�$7�&�wvH$d)�̍�^�^��U�b]��&�p+����b��j]�v_S�,��=������"�K+����H�{<�l�ȳ��2�GS|ɫG�E��ڦ�k�nP���YlL����c%��޻TO�2����U �������J&�x�q���4;;c'���m�U?0�	�?A/m,���
'����
&æF�^��K���,���I��˅9|�#ٰm՗xȉ�=�J\�4�V�h���)�u�|�o��q�0��W��K���ޕ?Ыҷ�v�5�թj�u� c�b�6��^��_6��>�떨he�/Q��u��20:��.؟�[���o��qx�T���uP�#vǯt�Urs�B��X�n������<|��g��V���z���jp����/�� ��"� �͉_�Z�����H\���=U)#P����~Y��>��ű��n.m��i������c~aP�>T~�����"&D$C	hM�gS-	��%WG;��t�z����<K��*����y��������~4ӿ�W0���\B9��u�Wv�JDH���.n%�f)Bq�pw5�+��[�!��I�^�/�v$�o�ؒ��	�&ؤ�lT�C�8-��^�{`f�v��p�\��i4�d��z���\�d�����rt0�:/s�����!nY�G~���OJ��@ Y���{���L,>�b4+�������X�%b���>1�rD����%Te�ٽ������{
445模��/�C��L��R<��,*��)�%�u�%p�%�b�����:����A�I knOxnv+W�ݠ�<��;		r���v�ZdLV'i}n;�e���V����[$�F��Jˎ�l�q��e�LH`E����b���W,�x'L��[Ak�xy:����Z��n�⋾��Wz��f*�!�f)��t�c�����ܫ*9ε�]gˤf25ă�c��h/mK�{<�{��'��9�Z��:�9�:^{�솿0�$'MCIi���G��|&�8s���b>����l�޿�4�*#XJ��0���\uF#��=�[.�ӼW����ٜ�_y���c!0	��:��&��C�f����4�_:�����R�Q�!/0|&~��j�^ �K\z(��Ԓ���E)9E�?~3���*QK�P�E�.�3�/�2��`8��-�#9E�Kz~�g�� iIڮ�f��-��Wb
�uS�vj�
�XkO�X'ݻ����?�#��	 ���2=NN>c�Ab���~�_i,qbRe�e"J;V��d�J���e�.�o���ުI��7S�c�h443)��r++�u��&�p�ґf�5fJ-
w��KCo�AA2���0���t,y�z��t~Mn�\��ӽ���g�E��LGW@��e��۴�	CM�Z4�����&��~i��.��4�3֦�����86�X,�=9/zC	�^��<���2U�O���i�Ğ �����IX�^��]������l���M�E�~�h����G�ZP�T�׬����L(X*H��mQr5w��J�P���\H4�7����1N����L4�\���k�F�0����:�s�W��,��k�?�f��J7�П�Td���D�0�'��^A��2����w?���n�t1x%�VѶ`V���~�ʕ�{،�TTUZ�ku��g����E_�2�Ӹ{�C*�+I}����J#��ϑ����ɇD�*a�wp�>��q;=+�6��PSU� �{��L��M�a��'6�[y�T)�.�}�%N����)��(���A�4���[zf|���໘�A��7M�$��*��:8���y�*�%���uXu�WOȻ81�%'C#�Z�m��u�����~�]�p��
.J�S,⳵�U҅<Cb2Q��������bn٣��Ɵ��:6�9i�3e�S'�CDYbM��S9S�����1���I��وG�&[�V+�B�?�����A��pgB�v�>�Gƴ�Q�BnΚ0p����E�2��I������X �1m������adG��	��i�!��~�f\Ԭ��w����g}	?~z��]�8r^q5"��S������H���+�}�)�K�g�ӯG��M�W�Y�
�L�~p�}�j�;�U���(�7�\�C`�->˾��w���ƻ�`��o�E�i[t��D���P��Q[�7ӭ�$R�T-�g"PDm��$0�Ǐ}�R|z��W,�'ф��%=�$�rZ���6�B�d�G�ezQ��n�҇�>ɚ1נ���A����x����&�3�1�ͮ�y�%���n��u�Fw͔�rt�3[GRɄ��Y?�@����ٓ0�}\�d&��j�S6:0y��/�]��6����l�;�E<DוM��s,�O��(3���v��<O�����<`��<��mv�\���f�D���,�2�]>������<'��>�gee�x?���8�D[�
�9	;ji �c�<t�B����lUJƚ�R�/����jg���͈MT�!<;g���/@�A�Ģ���<CKɕ�gz8�T�f��IP�}Mbؿa�s���|I%4��Ϧw��Կ-/ȳpGݷ�������s��x�3Kk>�LZ�Ҽ�x�r�@��^���t]J��{v���P������L�P���xX}L�VQ�c'���`�}������3�a��O�����o��'�ՑRJ~í�@L��`�!�(5�B����d(װ��%�H�Zs�ʩS�i�(zL�̲F8�6�$��^�3������LNP{�6)�\�X��P�wF����ȁ���|��d�`��H��2��7��@H����|��8nHПB�|�k���A��� �nl����o�X+�q�*��-lvy)�GJ-�
�l,�r�6�[���S���ZS�z��^!7ЪlO_�ӈ)t��A��/ʞ����_��|$�;j_�F���Րj!��k،CH�H�c�+�r���i�T��P�嫻�c}���
�>iY���Q.t�7�u|��b���#-cp�kTϠn�,������Ծ���I
@�<h����}��go�D�a���kk�d��w6����q�����6�U�+o�FWG�a�]��ۛ��b��0��[2���>	�[�T� Ŀ��?�D�k�YzMV����v�9M�����Bt�𲊊�o�y.l��9g��V��Bg����n�K�%����ӣKŽ"�#>od�����X&o��[�Ք�T�&4��X�8#����/�F\�Hiw��_Hv�>]���������dm��;:B��.����A(eE�_�Z�2���P��xQ���v9W�]Ffk�
�1ͅ3T���(R�O�]#}��n���)�k�-�w��YC\"AK����<_��m��T���xBʥ�ndH���O~d��8qt�Q7����n���[��w�u���X���e�l��zJC�W��V�de��[�=n&$�����msF�O�[-�8]'�碔:�j杍b�g/f��"�4�t�kBc&|0�Z�#NS\���3ӶN�!*�/�9%�ۅ��յ������U��u����Q�e��	����,+r�h%�Z|�L
����e��Z��_ؠ�JT�Ko}wI��7W���		�W��X�Qq��~��Bnd"���s+5�~�0AK�SO���e�!�Bc�'�����Q�#�F"�n�lo�U:Ϙ������H���?�y��q����t!lS�9
q�\N2�?�_YW��$������Z8�����[����^�A�!��~(�f�ؤ$�Ms�2�b�p5�-M�O���-h�Sud��9�-�HX�����+�f�ip���;����;���'Hz2l��ى�K�nݜ�!�3:fO-Fc W�DbZ߷��!�W�m�.{
�ʮMQ.gr����߸������G�;>�(�H��KMO�/����:w�Zg�W�����d��,`����;�ԏ-޽�?p���`�Ǽ�wGGd�c=�?G�G[���������\s��>N��sM�
�U��7S2Q�~hL����w-Ż|�'�^(�n��͢>���VnU�r�H�_0����Z���s�z��Y���HF��'��f�*!Pj��戹Q���B�<������:=��A���Mۘ��������1��Q�p�(W�d�?0)�N}Y7��3ڻh_�,�]1�w/�S�O�1�y+:񼴊�9�ش��.@�m��\*e]����m���.i��@T�}o�DUF莖Y6���vp�H�����B�f�kQ6p4K��ZD,ېm���&,g�<��}�FG���I�O�����[���;����<#t�c\����S�t��hm�:ky��^0W���H�$�ΣΎ�����@�*�������I9J��8,�V���Y(#�_��#�P��~�Qw�Wֽ�-�:�cYgh��h��Hpl���\L^y��B����n��>Ș��$��'��7�8�j't�A���zA�x^$����g6�@����i�e�I�^���q��]��ǫ:c����UI+jQ���m�t���B8�����R������z&y�Z�0�Cjd�V{g�?=��.�q�TkSX���~I�":��]�����4���lUn�v�����~��B�g�̕��5�57�Z�fF7���VTk�3�,tqK��ܸc�}��xS��>��n�}>��H{3�����J���k��Oh��]}��D�d�ݎ�<=D^����D��,�I����<9�<وQ�>U�j�\6n�I��[4����`j�t�O7�ձr�|��j������P�M���ۻ��7���I,��ׯwI��|����2�܎ưX�Kم�o55/��&�� P_�~tTқ�jl�^f_�>�>���ע����S��4~�p�uM�{�+MKP��z��0�>6����^ŷ��{O�&���ϮlQ[�ڹ��ͺ��h���{���%X����^Z�ܨ��SEc�Y����q�Vj���ՌC��/,1e�dD�˙[+U+ˌ�A�����3X���_�ZҤX7��CZo�nD>ŭNp4=��/��UE�� +o��5vr�ן��3�O|irE�nmgNj�.n�z��@��x��S�C������X��)VcΣ��k�mn�jЀi�R�]�T��+&|��h�d��������\u�B<���;�vǬ�LS�K����OhR��~%�u�����'��)���L�����OLd�Ĝ|�_\WB%(��О���.�殛'On�1�>d/~U���:�}��y���	��z���(+֔M7Kǀ���/=W{v)|f���l�&��!���g�Q�q��ɵ��w�5��h���2�0�qb�h�V;��[v���^�w�v�KS��3���	���60��=�$�O���I�w��b<�}�,k��S�L� yUv����#��� ��a/�wV�M��2�`cG:X+�_�������PF����v-��p��Ȼ�N�$N`�n��Q8�;�A������=��\������}�MCC���F��_L▨��β���E� ���!����㎎�Bk$�5��`_�kaaa����@J��ɫ�������`aU?�Z��/���IR�l�k������P��p��{�n���[Ωa������u?�\��G�Jbe���M�z(��*�˖���5��LqeB<�,��/+��٧����	�������L���8$������o��Oq,I�vFu�LB��<�ݲ�@�_e�I��a�U͑���wզ�{��S#��;�캎���>k��o�F������w}�(�>���11μ�8{���
{�e]F��7�ag��X�"ʋ��s?
����_cyn}/����N ��g�Iq�����/����5�^Bl��ޛ׭�b>�ǟ�p�p���U���dMLpQ��JA�=���C�2���U��9�>�$�ײ�ob @g�R6�n�w��,���Խu��v�:�����=#(����7��|e���
�o=���:��I���1�G�#]4cS�y���̀:����+��ѶV��*�rn��i�%�^�[ �AEW��	V��:&^]N�1���l��Xκ�FO��>�V�~�ա77K�Q�,��7���րs���G�����*����1��v��U}s�H����	u��S������RiG��j���$X��LÙ�wD9�s$�?�T�xSj�޺�	K��~�7vav�����~b#��nŌ�u��������K�!���6�׺V#9�o��e��0c�>���']�u���\{l���������B}Y�k�AS��B��F3�ޖ�\)��Ҏ݋[��i��Y�5��=-�G���'Gʯ�9�s�eB�c�FK�K?x��I[N9Z�o7T�d[y���͵*��]9h<�K!���	�?�fF~E�Tp��s�ظ��X���;U\��Sv�7�7��ه���;z(p�KSn�����<�/W�m!w�y?��J�ȼ��v�����<��0�=��������dGњBCㅫ�%=&���:<}R��$N����l0RQv��眿ˏ�^i]��R��t��^�4�]��3	�K��u��)��ąg��y����Q���X	ON�'�w�"�g�:��FWVƐ[����Xb�yQ��ҩ���j�KV��D�ڌ�΅ɭɆڙ�W��6�pZK.��ry�p[�[��*�eLT�n��np��*������µ^���?N��岒�!���%[
�����\�{yC�?��R����L���]��O�U%�Y����g6�.")�aU���m�^��K��F$�����p���������Mc"<O�ɸ��:{�9�*{��w�b�x��<�)╩�����!���(Og�<���aE��]�0JS����%oF�`��o8(Z|u��#ా��6�R�8�LMM��Y���[�mlX����['UoE�5\��=2�e3e���:1v��c�3:�����ks1IC̠�*�8�ޘP2�g�kФ���M�Ԑ��v�t�tRu8��Nlm�n������F����΢��N4#���B͵��~�!:�����f:h�2Qw��|�'������i9;�h[CI�����q��ӈl��}����M�z���H��*��u����H��brn���;�~�����+�̋(���<��4��Dy�qǎd�
��-�u�z;���'_����i%@I��p����T.E�Y_����#/|�G��+ꎫ�.zډ�N��-�-��'�#N�ǆ����}IWt᣸���*������[3ʃfd���«��iae��
t 9�|�	<���ã[��,<���.�.�5����7;�N�]"����<�N�?��V%:^�U��1a܇>�k�� cBr��3jnH����E(��]<�[�°.�J�o�Nxa�r�V�ت򆠡��߰��u��
x��[=�D�'��GGzt� ��>{���<���O8�-Ğٷ��Ϊ�yK�h�Cj��X��7;/n���(��x;L���  ).�kŬ��%[V7��͢q�@�Ѯ�R.�A���kllM��$>N֗�a�G�'��'�����������Rc�Q��)�; \[�l������zK�4�%>t�l]}U���l����5��b�=���H�t�E qg�Ýu��hc��6>ԏ>JD��o�X����8ʨ4�����[�*�D��\����\�B|ڿ+���)Gue���_��Ǘ��9���(g��d��#QW0E�@�{p���m����.e_�?�Ԯ�<̾׎	>*�c��aqy}��$vi���1
��0���V�ޝ�C��ЙO��s��]���LqIm�dۆ�UD�Tu�po�_��dF݄CY���%��{����������ki����Ķܛ�8���m��{V�3b�u�r�N�������zM��dz��$�͠��%JZ򺤅S�� \�m46lK�]���A���&�%��_\���e#�D�n���F���m�~��P�M�)�b1��������&J_���Dr�->oo1�<#.b�q� ���f�E��b�0e�8�\����;�Q*��%O�v�����aS�"o0D� j$s�/�}}B�����Y�	���_�ћ�Ï������}�D�PȐ�i�m�T}����&%4O�!B@�/�{�%�3�D�����
!��� ��0�xf�����	���J8�<�|����NA�+�ؚ��g����Ͻ�����:6�׀�mu�m�j�#�T���;_9�x�����P�-�jh�!����뒻�X�A����I#CY���]�%�B��1UJ4\Z�c���Ո8��"�$��sgy�_h�4��U�&��ϊ��|�P+�����͇\�F<�ے�?��EN�sQJu�t"d��d`�qsrОk������.}�.&�;�&�(*v;_����n�Ϡ��%!7���*3���F$�	ߏ]���29��?��B7��՟}۵�W>���������:�)��eYdy�'�G��Z�Q·������w���ƴZ])
�oݵ�Q�z�6t��oߘbۑ������O�ֿ$��l�-8�{_eo���vx|�(kM	��'�]�\0�ǍjL$%���]��T�cQ6NF����\+�w�-g�x�_r��`�fG��l��߆n�'dU&�a��ٽZciI�J���Jۂ�Ș>�]�C���t)^��sjs/��"M$�5�(Ux/ɱq\S+XELMP�n�|9m.�\����-�f�+ rw)7�z�;[Dd$tu�T�6�/��Wڇ�(��i0(X��|����/b�a�g�Ӥ�^����U�G���L:z��ç^�>���3k0����
�� ���%��F����!
M�?FЏ���+�/ɫE�ql�<��4�o� :�2n�W��H$\xX>T{���˼ǿ{`�>40����\�fD����HL��<��=�sz(���MK!�s���vaycK�f�.�据�S��
�{����hm��Hܺt��]Ϥɿa��@�(���Ӆf�Z���ǭ2n
j~�;#q�$���D�}<�{g]�"j�r?K�`�x�~8���"�\����
��bL������w�������x�L^l`����nc7��|/����>�\�܌�K/t�W���W2�x����ݬ2%P����1��&�P��˷-�cy���ê��&a��"�lO�Ѯr�m�Ye�-�HTR;̝����0�k��eC�|��҈�q��<��P��p�������a)����=�����\��5gW;��I�x��oPo{�|�U:?��I��=0��}�ECp�b��u�bɀ3�&Y���;��z�������xN���O����OpD<���P�|�9�I3+��4b���j�[��%�8#R��%�  C�,Qn*~�AvMM�RRU���^^2�u�9񎆄�	q��/j�#��EQ�o��:��SA~[��1�Tt\Z8�i�J�Ã�+jjs��Y{��c�W0�r�Z����oN�e�������h��k���/>>K��f!5*��k�`�PI������Ơ���u��C7=]o�O�C�l �B���^���lr�I%N��W,.k��kPRg�
����^O��㝈�3>X���q^�B�Ux�͘����U�>
�����h�k�z�k�Œ���S{q/�,�����a������:�1�AH�b�S���-��W�erNghNWn~ј����;�X�.;�r֐,gIr���O�Z+#`��!Vn�8م�fg2���������%e%���|oƋ;/��R&�X,�=E���r������$��<���s��{�'h�2g}<�����6 $��Oj>���:�������׆[��1�~�� �$��,ʪ���[���<���ݚR��:9�����m�'��r�8Y�HJ�ƾ�\n�q\�8�#k�Qh�֍D�.�BN�rX=E�$~��-]{�L:à8J���Nk�Ew�ID�%�0v��g��;�����J�lw!�M��#��� :�s���E�;�g�mW�5��뭜�|��kG��+s)H�+���<��:����*��p׋ڤ���h���%9�:?6A�Y�|!v��}��v��^=�����7��:@9h�Z#_��<%��Qg%��(�ԭ�*j�sP��o���o.��'8��'̷ߘ��0��e������-����V5���> *166��ge}�#,,�́���<y�9��z>�IȚ�m�9F  �J>_�M�TC�3�+��a�;[H�s@���7��e��T�r�P����/�����rU"�h^� ƭB�ؽ��簀����S�ɝ>w6�0���:�K*\o�e���>����2�	%�G0��ҍ�?t���Q&�N}����1L��Ŧ����T���ᆚ�L>����^?���2��_j��i�߫N>���/�N�x�uv�V�NA�g+��{]��� ����u7��3���t���I��&L���.��������`��/m-�a�%=�큡�8o�뵻�a���㑬�@י��&iiIh�^X���OVso44�%��M��2F^ |zrlp��"=���pJ
v[��N�t�0j��M��f�0����� �W�Ltv[�!���).�ɚ�n�	۴*��[�+"��v�1SI�L��ص�ʯ��&8-�S$���7_�6�t��Ӏ���Wy5^��\�2���*v7�/���?�h8��������byw���I�΂��v�	ֶ|̈́j���MYgb{u����U�~!%)��Y��t�y���� ��5�Ny�'݃qq���z�5P�4�4=�5	 SBئ��/��aEWF�_��i߂2tm���:7�sff�]�,|�����-cšt	X8~�����Cw?���QF8U����L��J��$����O:�-��e��4疤��У(�J���1�df��	�v0N}�,�VWp�|�ݢoi�@�iQ�8]F$��S�b���<����]�����dU)����1|�1ǤJdd�I��aУ�����M"��C��L�V��{�e�D����ƶ�Ł?�D�u# �#�w���Hۦ�û/��$��Ia�h��6}qN���+i���A���� ;=mqQC��+��~�Q.�S:��W���­n���%�1םlp�����C������q���" �齖81���/�(��Ay� �}��w�G�!QQK3��f�bͩo#��;��n�W�5na�<��l�>�{aռ^��8܌�'nXO����cN�/��w� י�h�)hc����$��Q�i�G.�1G�j����KS�]ryE���ۋ��m{h������+Jd���h���C�i}�G�ZR\��+�ܙ�+���r�9���r#0YC!&]��W˰?�K�]L8V#h4Cjˎ78��N���3�7�F��7�&M`�D�3x�&K5����O\�B|ef�|��qS{�5ccIeݙ;o�gbV�o��bŜ�3�!տ٩u�	��P'��y�ߪ���XO��;����
�<���Ӱ@��l��}����ON蠒Y9!"����4���r}���B��{%�<�Dֹ	q�����5�l����m��i�?}b�=u���ϡ16f[�艔7���1ۙ�ƙ�޺3�n�71}c��ڙp��* d3�{A�]N�w$�t��!~���=H�t@ۨx�����`Wr���{��z��8��8]����?����ȷ1s�
��V�VFk�[0<T�0I��*g�z+r2 ��I����%��4#�8N��\R�����K�Z��/D!�;f�$M�\P!!a�ЄT>�Ȃ���{Zg������z�m��ڌOO��-ʓ��*Ch�����=�[��Z�HN�'0�d1?k���F��;ߍ�ݕ�bv��SPF:�af���oYZ!@ȊJ�Y%Fά�v� ͤ�n����x���_< �kĵ�\���/�9V�Ky��o�z�����wOS������o��3�Vi�������'��������G c֬�+�sqW�к�D5��n�e݇��o9�7���\9:�������$���<�Nh��o���C�^���� o�x�݌r�Y���ַ�g��K;���s�,&i��i��L�D��=3�w�F;�ϔ]O[���>�!<f\/��'ػ���o͑tA�-��h�6��x�/[>�wvA}���ge�p'K$T)�C�,>oJY�K#a8g���h���e:o����]�����Ŕ��JT���8����H: �ڞV~ϛ�;p���n x���&G�����������"1}���Nv��Q�����kyt�4S��<c']���5nn�;�W/[df�����3��R��^���+��� �0�	(��E,qR��ٝ�pz�Ү�
pX;l��&�(s SG��� &�=�;��P�9�7�+�8���ªV_�VP0�2}ǙR��8����H����[E\*�l�l���_n�פ�A7%���㫞����g_}�]��1~�����	�� ��}�Xb!�&����NDo�����7��X����;�~��A����"^�mk��e�?�X�碌����98�By�?�b�g��1��s��v�6��a��-^rh ��>!�RF�"@�Tj\���. 6.ކ��S��a���i�@��DV���~��g/��n$��<P��y�q����}p�J�K��u�AE���VX(��"΂~1��1�yf�>HDAx���l�$Df�,*�%*Jk"��e2G���3�	5���1�����*��e�x�=�׻hD�74�ԇ�<�C��2�B�ԋ�@�]�M볁�4�In;q���t[w2 4@�(eF���>=@9^�,_�{��M߃�O���y�Ω2�C��W�s���5��~��
ķ>]�I!��	��a��D��V�t�R]%�Wh�`�'�AkD�l�#c⹻e�\NS��2�+Q�M�
wL�lB�γJX��Һ�[�)�@��R�Z�>�L]�U\F�fF(_��D�m��5�s�:u�qq�)l�5�9AR��#o�A�����tϸ������0�Ah���<̡��T�$B����/�%�煡��������'[ܰL	����	\Jy	��n+Q\�?��g]ol��[�Y)J�\�hF��d���	�g�mD'�G�{xٝ���vN��_J2�����\|0ש��ԓ�w�`ΐ��㞧�%�1�|�jm����@�_Ƹ �[��C$E{�=�57^//�R|6r�a2�ϋ+-
� ��F��	-���i����P�b;/��W��6��㹔#���:Ƀp9 ͒����0Fmf�ώ"􆈐1�̡�[n���e�5Q%��
��9�=x�e�.���IA��Ǳ܆uwK膣Ezd��a�w�l�={��YӍ��>L2�z�xl�|D��i����%,��kv�QG��t���n��J)����`��l�n8e�Ϻk�'|��ځG��|G^[Ա���L���އ��x���m4��(r�xU$��O��A���8'�ثD����k��?@҂Y_h<�!4�Ɨ]�/V�+g���>�4J���J�}�x�VPF8c���±zA��̋M��g�|d��d����~FiL��cA�j��%�@>c:�+��Fk�0{�,.�ֶi^� �(y����>p�sSx�=;;���yѿ3[+X�qo�Hql^�[o�gvGN�uM�/��f}���Is��F�*-S˟F�}�H�k{�}a��`"�d��OT����3��A�hy	O�;g��ZlS@�D��Q���;%bo�6ƞ��hg#E�U_��F�A�tH7�)
H)�).H��(]��t�t#���� -Ͳ�t.������;�2���>���|��y^N�:>�?�+�mi�|��eA>TߠT��~0??�̟�o�~�	��~�>�������d�;]���W=���w����Vɳ�zKs�_�F�,~"`S��u�kRA����4�5>���%	��_���~b9�+0_u4�:8�h!w\������c�졏��'�e]L?K\��5���vN[<�u��H���ʍ���{�gU�L���b�PD�#V�	�9j1�F�|���qv̛���u˪��Of��fQ-Q3�)����QJ�T�5�t�lR�]D�`qÝ_�Vۗ�O���,n��X4���u���	h���O&	:e����JZ�$al�}g�H�#iQ��@��3I�����F���&�7�lFq�	g�5j�Ky��1�&�z"����
Oz��^(x8�%� ����+�M���%lm�}��N��w�ҍtw����r�C�/�q��̖��Gs���`G�k�u�!)�V�z4�����j�%��+�д��f��/���j��K��w�����nj�l���ߴ�����+�W�x���2/�p�r|�=a�b��'��g�����*������d����o*�d���x����f�ec�
`0F@���]�_cZ�i����=<���$�	��>l+}����7}�u�퓍�U��(�.�OO؞����0ER/�`�0^G��,���Oz=!o�X1��r�z�g	��ڊ\�����*k��K/K���/�g8�����{�./O��O��`n�&M�ۃ�+W��ʬI����B�0� n��+�
ד�F���ʌ	*�~��3O�/�G�J	�1X�-�����A��nͼc�zXF�i�7�C2�/e�6���N���#�6ǸfS&�_9K2*���9��PU� ����pA	��oO��
�6wB7��xK���3�TjĊ#��0y�H#*�[����.�V��v]�x�>r�Ű�w,L%���G������*wh�QĜ��i`vl�ߛg�k$�=	o{�֝��eo&=�.�g&�Ұ�l�lﷵ(/���4��+O�0l�Rݥ��`��$S�V�<�LtҁtWJ!�f�9�o�������bf�u�&��kjK뉢�̡L/Z���0;��L��������+שmwZ�2���4xl�;)�8{e�'j ��ۣ�M���:=�.T�Ѐ��H��0�.��������1ܗ�L��ó�?�/�F;׍��J�iᗕ͠�M�
��-��J��	 � ��1J����ܢ��NJ%Ծ��4M��`!�>�>⨞u~қ�)��S���V@tt����:��'%%7촋F׷�F���}Q~@W��٠�lXǏ�A�Ȝ��j.�Q�'��y�����'%%a`t)���	RNz�1���?n�>��*v��b>��� �/��1������K���l���p}���r�MҪ��؛�-{�9�R��S��﬎��Xzׯ_�5]rH$r\��֜Q���v"--��2�Z���}P+n�&�=�U�bV�}ʫ��yN�7��zh3�O
�Z.�:��̗�Gmٔ=�D��o\c����3�4���18��;����o��?�`��>�>���B�s�(�]����ǃHܦN]$��R���	�!Ѓ�RD�G�/q5k��z�$�L��zj�3�5�t�%**ՠ�}�ֱ��8"˞�c�Joo���`8]r�E�� �v�e,t3B�sn���\Џfu��ҨX��9�0��>=q�Oc��7��/�(��j?r�������I`� 3L
��Sϱzܵ�>n�
 ���'ω~h�9K����$��yм���U�e^s	����,�b��u�+�G�Rn�<A�m+�F�V�3R2�9D�:��̇�������桁�\�G=#��R^jglKn���w`խ���+����w�^[y|�(�SU����������6�����+���er����7�.�&�m4�wu�5M�^� v�I�((��}�ޣ\���=n�)���-�L#�h�dۋG?\����4�4O������
�	�*s|Q����9��J��~:��^��ߟ�Z���$G�G��]��Z�.3�E�_`����O���,�PN$=��,��4P��y��u�K�~�;(�|m2��|!qT�!_	�gy{7�� �^:�1{`�J7!:��'��\T�zA��İ�����/�N��*�j!�&��xG栗RP��=�=#�aΣ�W	J�۫NT���Y�z���hr'/It�J���T�{����u��@j|�;��N��b��S��?�ң�?8��f0g��t���%�d�s�$*����ћU���B���٭��?����5���uӼ��ʀ��r���W�Ύ#9&��ݗ��]�ß(Te���^���qG�E`T�Ys�Ik�Pgp���B�L�rt`z�g�h༖������ך����3Skf�ד+�g�M:rHZ���l��'sxyw�5��< �d�&br��/���x�߈S��Ⱥ��Q�g����JK��CV�V��)��e�u*�҅�02�a�[0����c�n��hz�|(��@�9�/��^X0=��%���x������.a����m��UQ��&0��?�[�yy��� ����	fMϵ�ټ��<ݩ����]8�Z����������fD#���I؁�ɺ���8+nӆ7�X����α z����D��yL����L���ͪ��S���� ��������(2NAQ��#_,���Z1=e%��;�QPS�ۯo�@֤^���Sֆ�&l�(�+�O����hf�W1t�J�������SW��-�]����_4Н�a������"��/�;;Y�C��4��0CTf�-���-%��L����ϊ�`�.���I���G򀿖N�>V��gK&����4mx�x�j���.��5p�J�^�)帯�A�1Pm�?�	��QjP�֫���ο1�4x���|�?�d��&�V��cA�M�IR������)����f��ͫWM.	/)�<znӭH�uuuj��[x�����OA�WC���˽_ ���lf�bIX<�_~��
��������t�)�b�T7��ñG>�{~s7}�1��b����W(�+˿["8Iq��h���	j����n�����@M�/��c��9�*"}�/��jS~P�8�{���r��o��
�K��^���ٞv�K�Z�׎���(�����	$�ڟ��6�_$������	8��TZ�d��z,6Y蘿��	�#������kX�BЗ@��g����=_�0˩�p�KJB"y�/����D| �f���u�sj���t��s)�7��U(:�֪֡f��ww���M��l��?���U�>��R=�~x�zG��W��~�d�e�ե���s���6���y��p���d\=QB�_B�d#�L��3��]2m&�i;~��2Iqѭ˴�D$$p�����i�&UC3���.6��Z�!�હ���+�v~�X��o���O�N �P��K����$��&S�ne��25/�v�$�q��az��ʾ�d8eU /�iT<��bmt�%H�M�����Ә�p%oP���k�|�8���m����qS�4H��^��bLb�2��Tط�nX����?�u���z\�Pe��U�<�Ү}��DZ���C?v�*!��4̢t~j���E��O�?���2tG�F?f�T�avW&��\%��B6q_W�L_���B�ޢ���ۈo�vj��X���2
�u�x��g��ҵ�ǷL�C�sS������q����8��|	.�mX���}�D�u��Y���mʃ�K��[2�d��>���;z�J�����?7;�%�htf��y�j%����=Ce����E�0ڳ�clek|��J��b#�m��ҹ�����A��]��C�[��sD7��j��;�)H��^oMb�����Z��w�U�x��Ȅ�fP@`1;�L}��mp7�A�����:Qx�9~��i�8tvLH�˔���t�P�� ��)���Y�㍝�S��ț�N"Moӛw���ulm�"��>k�x��AgOlpr����I�;��u}�w!\*c���.�(~SV)1�����������t�O�V�a���`��8�����,9�+����z����sA"}K�n<pd}?���Rz��!�&�t���b������So�ĢP~���ë>$c��M[�R����=���k��'���G�`�bg�����\i����B���Dڂyn�R��2K�Ϗ��Vwn�����2b�a+�`uˮ�o�$H��������ӾR�ܱ�D���$��%��G<�R�fj-���X�-�RJm�H��{��8��XI�$qj)9�A�/�~+�(y\2Be��=��@�5O��J���/�9$wq`�{�-����^���0�vzv6�{{��+�I�[�rE	�y�s�Z�G7�z�$�[CXgwQ)��C�b���B�����P�u�%Fq�Ge����)��usV|�eCRB-n
Ov�ަ#���y'O�}��	]v����%a;CD>�S��[��3�RN�!	$�:����XR5�\vI\�t�/��*��A]��<��}��Ŭݞe@���_Cg��l����]m���Z��YA2�9:hZ�$g��R�47��5��(.�@�XtJ
~��m.���s龺ݹ��$5���\J�1�Ҽ#`����n�K�V�Mq"�X<�V�9�8��n��/D��6r?��J��gV8޶�V�T�z������"[lf,�'G�����U�����Խ%jo0k��@��hM�"��Na3��s�o�x����a���1�&�vv.05;{�	o��q�r���Xս�7aByF�\�W/�Z��vv�|�C�(K��ڸGts����Z����0�c����as�}]0g����	�{�@��KM��l���lr�1rx����6��e�r�JL.Ԯ!�PBϩUpxTi�?����_�*B1��_"^���~�2��fO� ��h�~�.�����8�쵺=���V�K�6Oe�%�e���(I�#���t�t�!)��"@W��oN�6��Do�/��J��o�B�,��W��gBKʘ2�Y��<O���/�̓�����Ѭ��� �_[�k|ef��;�o� E��]o��2r���^����y�߁z����kh�~W�}�LwG�݋ɞ�M����^D�9�M����k�_����~Ҏ#+w6�(1ѿ�]����+��d���Q��L�X<��Um�/
w[4(��CR�t�@L���f�.|o��VO�A�6K�IG%\���Df������ck��)_*����4�{���k?���j��NrЏC�%�o:��(�xH}��fX�:��I]�Z���sN޾�:�����������o�LDtW���r���;e控\�wk��X���l���w��l�����$-����v�;�J�BW��!4���H�S5��s~/���vg-(�^eċF@I�6�NfȞ�l�>�>�kd��9����z)�������JEOO�{C�y��ig�6¼���rglt�I�ުZ��n]E:\�3�<�j���6�s��W���I��M�qK�"����e90����W����c\LD��g}���H��=�`O���o����)f���96v�S�ۅ��%�>$��-~�?-5��1��E�$��ޡ�&�8��9���ou2<��U�lݔiH�����cz�=	�K���c���'��d'E�F+�WM7�0*iկt�I�[T3C*��~�	p1���s��v'�_�|�u�:�Y���u�B��T��T�k}���Q�O��:s�����
r��w��)�wf"�^E!�C|�&��B�J� .��.�}\X���tB1�៙��f��W�L��U���*wPki=*�3���q�i��)�rN`m"��3�$^3��X�d�����o��n���<�����x��,h>t���� MT`�W���0%gp|���Ԓ!F��}�ao� Z�^!�Zx�p��-�fM�U�E#(�����˦`����&)��沌�K4�h�,{~d�ϫGߍ������K�m�^NVA3>����D-����Sծ����'y���������([��88h3�h��`@lH�o�k�P�шG�@U�y���k2���U�D �lȓл3��,�!���������ZR�E�-z1�_NT��؎��De���,5�$�����z:�g�z8����į����G��j�'�tuu#�8B��p4G�f1m��ނb5oW���s:Sc�Fm�|�D��эT��^N�Laʣ��H�x��є7�u>eh`�j4� !T񋋨ܢ��%�������C_���)���jC�+�J��z��bk���H$>�wû�➸,Z�x���K.�lV��D�� j���W�BE�6~�e���Ncͧ���Ks8xj"�KՈ�w52�
x�&6���yl�P���ow^�I%X�#�h��ݨ��W�B?�͘m���pOPH��+6�����L�7��[n�Td��)��C�௦���3:���/}�Ĥ�^��!���,7�譀�E�e�#g�̯I���.���S��6���5�c�<K$��0mI9#u�����?C�ȶ�٣�B� �m�����\���Ob�wIȊ���L��+(�dw߱���1���ߝ������0�r�n/{N`��s��r�~afV!E|%0P�L���+�o+$���I}4�mv��9\�J5~jB�vk��q��;�?X���ᩒ9/�ð~H�7�((�6�6w�����W�'�s��	���Iț�?�7�B�T��8���o	}7yҏ�_�qR3 ފ��poC����sΤ1��E�x���8%d��T�Q�[B߈��tW��8e���	]����iS�I�� �Sv��U�Y�$��5��0?T�
I����^��UA��^B���K��׸��R��c��K46��Kw��4��`�+�
��'����튍�8���t��N�4Se{�0���&�^����8�ק\��EBe��0�����,��!����
Ǝ��\B!���&�!�X�4�zw���>�|��3ڬJ��H�-s���g�/���=��}Z1������|Qbb�]�k����ڡ��|���N#��+wr?�
�i�����`��$x@��!�mEg���1�,Q��f�1�dswY��.�an�'\�;b�,Sh�dG5FPL��v���0 ��H	WVV�Z���[5�p�L,L���Q\�'=YIH�����wk�kD�n�<����L�j���C�.ںl���ġ�UvP�Xp�s ˩���qB?��� Ōf���`����6��^S�oꪒ������h�P�\�鿼���;���f��
�s�����}���y�PyѪ�.y�������N�i�+�Mxk��w�<߯j3C<]<��O�p� ���A=��<��ތ12�(���W!����h<d��Ӽ��.�̭�g�?�Hgc҂�ؙ����d垝��K�sʬ����)�rf6!M?/��3|�g�w<쩤�"1Y�̨�!�������@P�ʱ�$��}das�2���Wפ�w�M?E˿ҿ�a:�4�ů�/��L,�����G+�-7�@/�~2�ؒS>�Ǧ������;c�=��Lݓ�. ��"�ܦh�J�A�d}-͔�ʔ�k�yF_�l��DRٺ�G�3������1#vc�� �8��^�6=��8m�.A
�4oY9-����q�_���l~��:���k�� �1�_i�|�/.���"��Ռ�?�c�}���p������_O�x����!�6K��5wqQ�5��<���/)���2$%L+��������ء���L���RM�޸��g)����?>zA����������r��m��KL�c�&<��s)`݆���.��r���6mI	5i�D��4�_���o��x	�bO��ʯ�av��T �	?`�c�?�$K����KD�ۇ�a=���yRm9�7�i,���n��oO7�j��Y-gH�o)K��D&�q����#P�f�?��L���Q����C���}�7��$\��ր�ш���S���,���J��oʸ$�g3�ŏeԌ���}��Ny�����/h�HiU]ޥ�W�Na���`պ��o�3�2���]l�/�6"���V��D����o��z�����Ï'��<�)4l�
n��{H���Ҳ�+nm�^I�?����<>R���}N �
xǧ]e{'в�U�z��ן)M���+kt*�
#�5����� I# *��:�L�m��#��(����)jH��z܆R12�D�-��y Udx�cI�� ���6ZA7�s��\����/�!�p�=Mf+�9h0[2��-��u8�y �AbT>G����Fx!(㾡ߠ�`#`��[�)1�p���̦���-o�ct§`O��YT`��GTM��C棞|�򋷵�0pQ*`t&�65�T�w��I����9��B�����I
=U�;6x3O)�v�����cD&���כ�ұ���5���r�z��l7��s/3�r�J��0�<������������"TC�"'�p6�f����(z�q��m�N�;�-���/�a��W�����I��t�pf�HQh'��*�2��%���"f���;���������q��J�	`,WJG#����RO"s4���"�/H��Yl���8�������("�KbY�{�ۛi����a�����]�|ӆ���ndd��~'�!��D�ˌU[��ޔ�8���8��Z64d]���fH��S�D�����J1P$�`u��5��H ��F" RS9���IQ��.�Q�砬�2�:B��-�ȃ�s���ܾ�K���T��x���+Aw6᲍ݭΘ�!@Ʒ����"Z�}�rM�@�]Z��Y2h���٩A���O<���!�S�d�Ƕ4y��##8g���<j~�f7S������C���5X�Ϟ�Ȳ�ʝ�g ��&w�����N�5�X���lܯv��X0��M��-9�}yԫ���&ɦ���T&Џ���x�î6�	��hۼz��\��T�#"�xҭK���M�gI��p�Ͽ��9��Q++��B!�"��M���|�b��h�*O�J��f��ު}}u��Y�@�M�!##P��]�b@�um���O���DT�FKG��*�VH��|�L�=�نm),:�5l�E.�L�7!��v�������vM�ߩ�c�S@ޜ���-,:�MQ"B$���@�jo����DG� C}��Ϟ=s��.Y�t�ś��ݑ���e��;�O�x~���K��y�x��~"�30�k�e�[�$���(�_�--M*�pH�����e烏7 6�����,v9G\�{H
tJJ�D`�"�W�ؙ����Եy$�;�&=���B���A1���CNa[��"�s��u��}l��2�,�C߻<ȁ�����|�s�>���B�_Bߛ��W�BNr{��Kn��v�zV��`�@�$Ӟ|���90�j�&��F9x�[�D
'I�S��|RS~��N�;p�>kǳ���fj�����lѧy��vl���
��q�G��|m����ǂ��̬%�t0o���۸P�<������p���MyQ�p�^��V��M����pKy��'M1��A��������صq�٘���Om�ޚ���?��b%K��ӆ�U+�d��O���Y������Ŧb3D��L�����FT�3W)���̮o<��c�
���|�K�lh�`����FF���|��26��L˛���'�$P���CRrZ���5�<$��l����^
� >j������
�@FMV�������f##����oU}�?c��˪w��о�A�s鐮4�����BI����F@+��T�z	1Q�>�U��o���z֒����Q߬�iC6�m��(NvT�� ��U����ɴ9�����H�k��W�I��^���8,��m��}X0��F�MNB� &=-�����d�󬏪�yϛ�5����������
NQg��ɰja�`���:��f��,f�̀!�Q�-�q)�'fJ�4o��	�-[���Yb�O �T}o/ i���Ч2���ÞH ��^�o�f5��� ^B̩dҧ�w�^Ǯ��������
��`���!B_B����.x?_��Ĺ��_�'i�_�����Ʃ
v?��]����������q�o3|H��P��2$�|��[kl�iQ9�,�������&J�@U��w̌�Nn��un�-����[<�����x��^'8�����I6��"��V������`6$��0�������G����U��3Q��x&�}B����ǂ�� JbXV=)�i�/F�[��8��7#�cF[e�==@iՁ����u�/z��M�6�PH C�C��p��~{�g�n�`C*�s���$5����͕�`��T�M�wm��Kv���)B��٦ |�$ގŮ�"�S��N&[�:�?_驺g���H��
rssf�YL�ͧhYA&{��+aǊ7�������e��-? ���M!����"�r{f��A�������r�	�"���6CZW�o�7f�!�Owf�)/hz�gQ(�r��{;	@����}Q��8�)-+C �5�*��z��iK E~>(8R�r��3�'����|��M�6�T@���1m2���R��.Z^"*����N��IT���y
*e�\����K2�u������/�4�*�����j|�}M��n��6��Y1T
ȯFR��	~y�a�x+��裢/��biUl?�E��������)�uo[�����Gm"�˟M��O,VV��;z�؏�b?���&�l��^�'
�'{\>�6�f�H8��&�}������F$-�,�	ȏ�����]�S��;�Q�,�.����� bLj�&�۽���L���1"���T���2��0���.���TS���s
��;8���sC��4G]���L�[����ҭ%?�խ�ݩ�h`(
��w>�f��	��TÓ��[ǭ���'{��8��dP�55��C���<���� ����U�Rs¬�ͻ��/FEBI�r�_����P�~�H[#�*&�y��^�{H��6 ~{�{�%�s:V
xN.���߭�X-g�醍N��iܪ�g�T㕁�;��h��xG ��[�UW.}H���߁ر�IϳۢӾ�������ls���V������"�Ņ;&�+OƏZ�o�I/��<�ř��G�r�j)�S�GP~��d��~f֋߂�~c� x|~yy?=�ݭ���-,(�����	�3�2���KVD���.J�����Ӓ����V�l�;�H��1�Y"
+��Yj��OX���uu�B���b�t�����!ֿ[/��Ҟղ=�'�3�>9�0�$�pf�P~_u�T�����񛚇c�N����9��<mQ}��1E�&�V���uboM��gk�-*kg����MQ�� x\sPfq%��ۦg�,L`f�V$g�&�ܴ$��cg�KcQ辪ݒ�C�����}��<�0M�@����v�F�-W&��sc�A�M�����vo���4�@�S"���ʝ�����۟Ar k�2�`?%��.����Y\f�mDLazd~�َ�w��hF���F<�]�)�O͡������Q�Qp�Ic��wnY�w�W#���gC~ȟb$������4݄�0=T2��f��:gb]�h���_h�/yJx�1}�ʹV�(\��7i׾���ѥ����/-/))iW1[*)�4:���Sĵ��ig���N⓸����������}��G&"�+s(Sq��:���`�����]5q,֥���B�i+ݟ�~���)�߮�M"�koW�t��dsT�KF �	�lc���w�"A�����ˏ1��}�Ɇ��z�-��h�!�Ϗ�"���y����A��H�ڏ&gC������F�v�n/�5��W�69.�ǯ�oQY�.B�[q\?�P+d6�)굿����-�;���v��bs1���'X��-�<�,v�������)�g�Y�H�Q����4�B����蝧���6=��O���}��?�O~�a2�WPX&��'C^�S�b����VU�ʏ�+�"yg������2�K�Yg�z
:aP�"����_m?ا2b�r�'(�R���*�f�r'�f>[HPP�X�Ր�����qR�������r��J�Np  �O�#�B2�AQC�S�����P�ϖ[��s��URҜ&x>���}b�gsl�'r�7�y�Ec�IM4*wt����p���kE�G����"y��\B۹60?XK'��t�H�����ة��B,"���	�^�dcB۴U�Gh�+Iw����,������g���l4���a���MQU��-���Q��f�_�~�)�0�䵴�]<؆�g�ZRߎPK��Þf�4u ���Y�\z t��(�g����c	�91e;�x8j����ڭ���.?`[\�(=J��rRy ��q�^j��F*Δ�@J$��rՙ�+�
�Z��ׂ(ORH���-q��+��w:�l�D���D�~���층���0�`]�J�i�VG6�Y�Q�}#[ku��FR���wT|yy�e���A���=>��=tc���[-����~����˦�"5�����G����T��)ξ~~�W�*�ff����aJ+6�����:%�:%_?��z����=oiKPT�M�����o��XN�˓�A5<�u�Jj����E���,''7���}��}f!y��Ԟ���K�'�O23��1��?\�/���Zj��kp�ڥ�b��r�PJ/���p���ۗ,����#	=�f��d����^���!�����-S��j���O�@����>����s9��%�kF֚�f�L����[�d�PlE(���v=t���B� �����i{��s�0�zEG<郮V�Ov�#�Z�6%�פ�7Cm���1��
�ϩ�?0��/3��T�n��=U��>y'-d׼Y�*Ruj*�A������cM�����b�WɈ�( �$T56q��&'�/d���c
W�uzcO��Ч�K���Upb�ׯL�ϹȠw,,���\�5֐Xܠh�&Ƨg�В#�77�D&�9����_ۯ�
���1�{^���e�T�B�o,C���빼�#]Mc����D��"EϮ�~�6�vXPN��
� �����OGp<�����*X���(�r�\��,��¨�s_�����R����k땯���ŗ�KKK�����U��V�����C�M�66�w�?�u���z<�e�{�-b�w��G�uuq����匎��g+Lͼg7��I���A�%�1��	b����2q^n���T.��R3���K�-ǎ�����L]ZZ��:��?���=$@s��!�pe��kcG�]D?���1���6��9�˝��������I����ЫgILc�h=�A�>����1n� ���h˵g_qZf���/��F<��M�>*Z��eq�3)`ڝ�M�@���ƹ����:���;��|?���[R��Å�e�����,x-N���'��k��Q�M;�i�gҧ�>a�HABB�����]�Ԕ�뗠�guC)J�;?�X	G���/ܜ�<��d�+��:Y�R�z�6����p��������4E:%\��x��  f��s�gk��;z� C�*#.��/�]Er1kBi��!�o�&��[���ʅ�I�k�Z�x�̃a~��	���a�2�d�,�Mj�b7�����d�@��O	�����e �F"���V1\��=N��o�bz�E�/�J��{��D$ͧ;ס�/�Q*ϞˋF:î�n�.�b��c���*�������/΋�D�T�%.�uי�[^� \�w�4�q�+/�i���`f��/�49��Na�D�!5��b�&<���,�mHe~m)̀��ڿ�½3����'�wƖe {e˅��ݹ�G�FMԀ�{�7��	ikV��*G���j���b���SE8��e�>�A�uK��5�4Z>m{HϠ ��4�Wċ�5����	9�J�`+�����P��B=�0867���N�[�P�^�
vo��3f�L�5]%i��)���m>^HT4��p����47w��@��C5^?P�^��ş㶢:|c�3�O'M²[?-���g��o}}}	ZE��9��NP�dSII	�Q:�ysl�p�h�H����$����BM05(J�FT�319L�"��Q��>^U:���	N֐q�0e��ƚ�6�E��K/�:�a�xF��@R���3̝��a�X���H��'����L�s�=��⦸IE51)�.��p���ƷC����<��q�E+�eJ+���p�}y i��=�M�.��uN�3�9�r9?�?��rT��SЩU�"Z頳(;�F�*\�j��<߸�=���q�|w~�G~s��8��5ݿs��1Y��㞄dǑ]�6i8M�E�?��2��ňw��v�4�9�S�9�>���)H j+�"�GMO��Y�0�`�h����~�^;ȏ�ZWz��M�Ǿ�Lj�^��(뾤��Ѭ��*G��	�L����m��#t������+Td���Y�Y8�8V��ER�`lQI�4�g�7��!6C�f�o�j@�Xח���
���W��b��XϓO�`G0�b�t�a��e�.DMٳAĜr�+++�'�8�
����O�%�h N�:�F�?IO�%OP�b��j�
ʪ�x?;*���I�j��� ��W�D2���Kdzy4���!�)��IŬq���1�r���� kq���,f�љp���u{۟)Y>����oB����{B��^��[ �A�w��v==�o���ill��*���H-�W�@���8[� �]���F&�r������#�2�+<�S��_�4�Fv���4`�6�t
�j!��9���#�{��_��+a��.��X.�~ᴸ*�������3ҩ�e�pi��=�,�x��B��ژA�ej��2N�_i�(��R��M��1P��㸉��r�=�r��� ���ݮgn�M�YJY�6*d�mK��[��'���;Y��4?�����<��LK:�s@g��il('?�*.¦���6���7kw�BJ��Y�����݆͔gw44�M�0�&R?55�>���p��6�dQP=��e�g��%�&E&7WCX__���O�%UU��L�΍/�FZ�*���?�����W�@�g��t0�ǭϷG�x"��l��.+ߘ��G�ES��(�;ȝ^<����LO���'*�~�Y[����%x<kb���ic�՗��c�fy:dmL�.��)��x�b͕�߿���o��:~�B�z��3��%�_0�'(D��)�
6b<u�Zm�)��,ە��nk[/�9�c�[4��E��i��JOX������s���5���ڤ�4�Q��� � |X\�no!1�s^�C�w���'-�C��k�>�l������pձ��m��R��~b`<����Xud͵��W�i0���L��5Ng����5�E=?�h�V�5�ޱC��W/�,�~7��$�U~\ss>��$QO�|1*�x��2�JD�J2����]�XW���}�͔�'dz���Q��g�Ⓠ���]�fл+JyK���N�&�c�b{?s��\L����w�s�^H��I���p�T��������V�~(��խM���s�4����m�`�y-���P������^#�[/��m �%矁�=2l�lp���'-y�x���w���]/�Fm��w�% ,N�;�Ⱥ�ե�'>����>�=�z���߶�xk]������s�����(K#�H�Ji/uj&u��]�P�dEW0&�ߙ��B�pz'��|7���?��U%Z!:��Ѭ*q�:ؽ/J03�_"��
Z��Y�2��<iA��)&��ڛ��iO����o�,R�q�t�cv"X'��ɴP�py�����I{��g5U/�elT�2<�b2��������0��ppC���v�t4+«���LsG�FU�.�A��q��*kj>���M����3 �F��#ej/TU�[=���z��e�N%���G������RS�DZ g�7a��{!|��p�R�޺�	� ƽi����1���}{[��&�$���pJ��B���C2FG�M�F\��.<��6�rlR�P����\ �����6-�~��VQ�'��O��&�0�,R��Y$�.� ��Q�����	|Y�Ђ5/�x�YB#,���q�MD��Gإ5�t�+}���P���i�������ƕ�uz ��q)
�o{���5�c��qf�n�TgQ�4k+� ��׍��Я"�w�ъ�[�iŤmt��ۅ��B����	tQ�y��!��g� N�U��EY׈� 4qȩ�_�Q��;�ׯ��y���'��ǫ�X�Ť�]�p�;��K&I�;N��ޮ��ωK��o߅�H̶�9��ɛ�F���D�oW]^�O��TEj��,C�?	֌��z�t{��F^6@u��b�jH�H�-���~�pK
����
=6&r{,&�i�X��tꦌ��5l[�,�U�9������v�, �l��K�B;ś1�u�l���MgVzU��W�"x�o����Svе��,�����ͽ�{��&p����2U�C���XO��A�������چQBR��Q��NA�Aah��SJ�N钆A:��.)��n���������pf]�>c���M�5�*Ua�~�p��2#�wJ6��1��,:1�$����
����j�i�}ϣ�A{�n8!��x�J�ۿC���)�CTXXX�v(QktD����腩l~�}�����d�d�Q�:���U
��?���\��e��74��kqc���DFm��a�~��A��",�
P�b�p����/,��k
��\��ٮ- ˲��|�.���2��sV9��|�(�Ӌz�nd�Z�ۤO�c#}/��'���^������f"m���hd��V��s C�}C���sD��)�$<�=�>l�7��(�1~�8~�ȝ��\���ƀˠ�ͫ?q������S�z� tt�!B��2���&Y��Z�������z������G�#F�E,�3n�xe)�w�Yۄ �)��]�B
(LC�����L����I��e��F�+�'�xiv����OmZ��C]����`�v�G�\_v��a�y)��{~O��H�	F^��KS���/]G�l3ª M��%�^���ῥ�n_�Ev���pw�?T���N1�2HǨWR�gv��z�A2��W�bM�$j�~����n��n>�b]�`�a@~��`o���l^ e|a�?D ��Y��1�`��N�8�n� �o��/1v>�Q��.� �>�_�?D�rQ��H;�cK���i*x��G�C�O��7$����j�����6
��(?��\ ���bo�&+"� lD�G��\���֣f��;Q�N��v+H��ijc���$��K��S<;D�>V�����R^�Ƥ ���5��(�p	�����(��ܕS����,6}k������?1%�9��j:�t`2��h���!×��:vuۚ�E��Nc^#q��P����Q#����;��B�_}cn.B��V}��A�
�%�77�l��Ǒ��|��.߾���"����������>-�ã:}�#��x����HrWG�B322�N@	�^�H�\.9��\I�^%~	�0-T�(l����d����8�?�KlőD���[��d��ϼ� ��������Y]�}6���O���D��u3i�`_�j�vM�?)�HHͣ5ƿ�,+32(���3p_��ӊ��V�O�%�+����ܡ������ I^	�(@+�%�;K�K#~�}����9Gʧ\�b5������-eaX��^J�wP���9�鮀=ےW����S��~q�/���킼�CAV�^w$����Mwg\�:��g����'�i�]}��#?m�s��']�N^:Bۘ�5.�w=�7�� U��X�������"|�QbW�.�׼���wp��4<<�1����I���&�
?7�"����U"�U�t��́�p|bj:T��A<)Sx�Y��c/�4��Y�.]屫Ӹ㵐��G�X�s�]5��'�`����wz��},��n�|)#D#��J�%�ġ�X���������>R�W�N�Y^!ۭ�U�b�z��H*��s}�O��i��[^����k����s2r����p���*U6d�����g��ݎ�_�W;6̴,�J��h�zNj��y���&>����`�u���!wiZ����f�߳1�i��اy�\��4����))K�����:	�K���kR.�@�>�����js���K>����x�JD�"���R�����M"����!u!�����^� #�����l��2���Kp�Q��mX��;)��xn{:�����Z�%W�B�	<�����}��?�1<O뚂�bk�&p�@���/��eCJ#�]*��<�A��p�P���Р�!��ɰŕY��M*K0�W"��7#c2:�l��ڬ�6�}C�OX���^�.'��ه\��5:��CbJ9)L*|}}b��h�C���j�N�R,����y�^���e��ʆ�c��k�9�X	 M|g��
nu���y�����A�?l�Q�^��\Y2u������=6��ʑXܑE������vw}3[G���U���\�ZR\�9�j��Ď��_����`v�do�h�NV��:P\\R�Yri��~�V8,�Xh�7H�T/�w���د��(l)a�h�Q�s!:k�-�fe�A��yV��
�B�))����9� s���H&Qթ��3M��g�B��/�R���Xt������!�j�d"��	�N2S|b{<����&{c\j*3���ij8@���	�A��TP��r��$���Ez7w�N��+�6�9+�TP�7`�x���ޅ�U�#uvv6�R��U�^���ڲ�aV���q�������O�L�
����&����Y��;dz�����O�(&��Imgn��Nt�C	q;Ġ���xmt;70�ۖ�D|�)�|�d+�;��c�75mk����[[X	���с<in|!S�k��;{�}�|k��h�aq��\�PrU����Q#BG3��3Mʞ�"2p�J�j��L�%OS�uJ�c����vb�E}8�:����4G��22н�I8i7���R�57GS-V퇅�C5����+�Lcޝ1���jG������海Eb�^���|��(�*�Qu��E?+c���y�u>Ͱ���ߐ�ޒv��sVF��E);�v��*���.���p>H^7l����t/+!zD�G�l}���Q�2>
��a�cz�oKf�-���N޶��׽j���.��z�����a����m�or�\��LyB�VP!��ۿnF%Ir�/�����;���C2%.���\s�ejCq�޳9�j�3����-��B8;`y/�>��6�M�T���������蠹{I�+}����J�CԊd::�KS�,r�WQm��lgY�k�;h(7\�}�ޏ*�3j�M���8�8���$�i���,:j��Y;<j�2K�KB�"?8��xHR.�,�(���yO,�h�+�����g=}*E��\�rA �	���_j/�Ş����QS�j�5b�]���4��/}7��>V�p_s��D���2��4�@}!I|� �Q#ǱUR��_]g��=�E�&.�v��$�=�׷�������.�il|e��y	�b.����u�D�N��9��x�6vϯ�4���rrr�RR��N��c��T༛@>��0?S�>܈'�)���p���V��̜5���:��켏K��
�"mU�Ǒs�avz��f���=��=?�낣W���6$�E�孛ە�K�ҳ&�N��z�\�&�.�:���}��T��)��-�iN����#�|A����k�N+Z��3���ǰ���;.S���G�8��$����q�6<��L�[����p�t2�>��|rQQ�S77�)g����T��c����4K�ٔP�	4��4L�as�+#�@�К���r+����7�D| 5����6]�r�SZ��)�M�l<=u���68��6ihZ���[�:x�O��ZB.a>�Ɍ!x�ū�UF�?�Wχ+Y�z|q'.�u<(z�्MJJ*�v)�n[辤�xȬVX002��ly5�w�u �,j���'ʴ��I���� ��_<��^��&�sY8&�K6�S
����ċ���l��I8m-�$*�n�!�@��-���
L�����"�_�fM������P���.�/��D�AP�E8�);e���!D��5�9�n����7�Qÿ��F��8A��\w��k��Ri��#����Ś��)[�B�T+Q\&Sab+壼��e��ι�n���w�B���v��s�ۿv+}����?Џ@,�WF��}3�b<��ϛlq����6��8��g�$��Qj�h2r��Q�Y�P!�BXճ" j%�XG��8*�� r�̂[���j8����}��W��P�{�P��ޖ2`�A�7��L<�o���I�,��w�aN7a�v�7�˝=g���(Uݶ�����y=ޤ�7h(y�MF�$�Fx�Q7�z0q�Cq$��5�w�&��4<�J������]�b��3�#�]i�ۡ���Ն�G�/`������(��3Ieī���<���^��q��h�\ӭ��/���+����_{}��2��)��}C��E��ݍ��0_Z�a�4��y�\Y�X����L�N�UTT����V�'rx�Ƽ�O��!u�	�<�
B%Ǘ���>�kǒzt�� ʧ��IbX;`NZ �ą��MɅ{����2-�GU��g>��ʒ#�(�]Y}�.����L�%$sPS
�|p�ԐD� �M�e���/���ĂJⳀ;S'�>�9�� �P��}���ǵsm� 'ܕ/�+%��3�+۔41jy�O-�7$e�N����y���%�E�S�g���C�	�����@3tA�}��͍6͞�|����A�~$F���(:T�d�e�L|��M����	m��i�^��?��ݹSGQ�!S��g3�:������X���.hO�o�p�[c1سu����WL\�8Yʢ���b�?�	ND�Ql>�:jX��
q��?���%����#�W)���W^�i�w�P�WZ
�d�5���J|�ŭ�QB�� .~8	���A���6��D�M�Zc�ޔ�Lx�vґ�6S�&�_0F�+1d4�q����,�	u�P��}��� ��5-M�6m�7Lk��1%,b�w�'���3���zF�^��L���&V?��ץ�ｦ����=4��m��N���I�����g�������ܐ��UF8z�-���V�E�Xi�	IU[��M��;;�5F��۞��QĶ���ok}��������.�b{�,9����{�v���,�%�Dh�^��ib����CӸ�3������$ciy�6���P*����O��t�[\��������<(���D��m������h�ֹvy ���<�Se�594�4X���C�Dͤ���,�)HT���Iw���}`5Q�?�=B�U	j|�/f���^��q�A�Sl��p7+�_�4;-id٬)G�
"}�A+<{� ~��as^�������8��ͅo��6ܦ�c��G��BW��7�}�J�_J��8o�+ ��,��r0[.P�t��Γ���v�J��(�S��PoZ��"�F�Ϟ��\-�w5��E���F�C�� �':��A������W+&�i����F�bO7L3���*����i��,����>�޽�s��UZ��I�n��[j�ZS�CU�H�	nR�����(X�/��X�k�f!��j��m}R{~�Ph����2�,ږ�!��PvU�*�OG�*Q1l��s�N+�I�������r�$g\h�sYVq�?�@qb�aA�D��ʝcn�|�f�W[�gV$$!]������V�{�Uqw�����]���w�!�c� ����p}�Zlw��锠\� ,hN��4Zt���V�n�'�W�}�	�U�-j����o�t9�1!3X@�
#a��1ٖ�;]�Š�b,�u��z�/�Ď�fA�?~���˽�O_�9f/"�0!zC�C�����j�X�`��O��ڇ��u�,w�]2���j�a�����<:��Yu�ygNa����),���FcxW���{+����jl^�xk�2��ޚ���@�U�umi5
E�gQ>�K���uH4:̯}�-�>�S�m��r���@E���C�zuj�:q�\܉MLA·�9�j��\�=1)���V�
"��<��«K=������L�g#��10��ph9'�.F(�@u4 Fh��Ghhe?Q6��<�����y8�T�5�`�o�|�/Rd�������hz����{������o�+?�a��RBF� �$�k����j%�w�"?�� J4)w���ͥ������g8��l��k�S
'� ��^���W����}O�'��~X7a.5����������脓(��P�Hdhoω�_.�7!0�D�w�jWB��kB���F�ӱ)�����xyq�Ț��<~�Jo��
��	�8G��<�9��oT���7�����:�YC~SD� �����B����m������Lۘ�_�x�@u���Ńm,�˻���!��s��LV����j�c�o��P�cC��`����W�V���n�y�����@��ނ�8%�Q��l�U��j�E�Ǜ�	á�i7�2k//��p������7Y������^��iȲy��Џ��t��:U���}����H(�n=n¿ ���]S�:�%��0>4�/���7i�Wx�TR��뭾�x��K�"���f#
v��_3<Ű������H�!)s���Y\Z���dڀ�|x��y쐼?zz�b�%e[���0�ipg=�����W|�:)魤��M�vl{&5�֡�G�*ax��&�(p�ٓܨ��6��-��/O����N�e��x ���vJ	��{�5���q���"d�æ�mh����k���}�G�������uE5+�Ϯ@N��ЙF�?�8���SA2�X��ɘ6�|�7�Z��!6���g��j~:~f�޸>׵�j�FΏ_�Gӵ�6�r�@<������b��\׾�������R��" P���8<'.���0yC[<��:n�B�/��O�zc�1f;\E�aq�|DrP���j��*DϏ�s��.#L�~DF�;�+]�����j��פd� �3n�ՅøLos?l5�C��5���hnM  ��-�t�oG�x4פ���=^PR=��H�/S�3z�!��*�޴�����;#-�A����^���Ō����\|��¤����`�P��`0�ө�����~�@��3�I#��<�7'��jAɹ��a�d�]z`��� �+a�و���OC�#���vy��fV,w�e�%(i����&*���rz��:C�h'�12r傿�{@�����XJ�~�Vd�h��4#�j��iW�s`VCN[H�K�{<��\��Q��TfV��]�m^��όc��lF�!�9ل NF�5��ԧU��~/Q��������ʱҴ�.��|Rz���5z1�k�����'Y�7o�"�R=�����|_�4��^�+�!i2\��I�����p.9fW�&ط����DOb>��ǓXq�zzH�&��	4x�d������1e�K@M<�E�p�x2utgw�;Ԕ��/�x�5���Cq�{q��`6%^�(�2̜.[���t�ƴ��էO�+��,ر"�b��U����fy������6E�O�����[�9�8����~��}!)��$�M~���hnc�q�v�L4�����p����q�D����Nh�1Ud`ꯧ[py��6Z�� s���m�J������=�����>����6�ΛՃxOˎ�t�+������ҫ�#��ڠ�Ј��w��x<d�DHn��i��g��o+g��m9b���nm���4�����Q,�iba�\�SV	寰��Jb���0���e�zx�+����"8"�M7�5�����s�W6C˽���%P��Ύ��|�9ʸ�����T/����E��=��`�6Ϭ9�
�8 {`��_dAA��Ke���;F��,Ow˅ee�lӯ���I�{v�fFSK+�ʁx�d`�z��}�LM��~�So}���]�l�\�p��C�gW��?�_m�0�}�y舌~�pZ�@������^�^����T�4C�:[P�e�ih��M���݁f�M�ZZ&��X�k]wdQ;����d��4Ѣ��}�͝�ͷF@N���������J�u�l``g҉�ߥ��Pbv������z�� Ը�Y^��Ϋ+��_=���~|{žv�3N�C+�Fڂ�����Q���Ғ��"̎��-n���9�|x���|��H������3x��n�-��*�����T���i���_��D-��w���{5F�=4�4��ض���kT���������Y�6-fU5��9��ן�=o��d�u�4F�!Л~�kH���O����m>�p��-8+��\dl/ʔ�J�~�o/���CԟZm�s�_<�1��0��yZEM^��:�c? �����K�I!�u��#���LRix)��qI��*x��j�T���O^������ȏ���)��u�~u�i����v�d�f[zQ0���q3��v傄"�d��Y��<.���qR�|A[F^7b�?~�D���{�l.7e����t~�?[=�H�O�)�.��,���r?8��^t�p?��;V�{/�4s!`BѰ�j���V"�U��GbQ���k�%o�Y���B�}%a�O7q��Y38�ٗ�qv	\�v������f0�{���ЋY���<�D�b�>GJ�6�������������S<�F*�"��ݝh_�-�x���x����a�5�h��"��`n�Mr�'�MV�c/���^��@��)�6 {Xx��^I�On=6ru���;lY�l}� \�)y����K����<w���)�s�ۘ�-�������}�A�yۢ/���ꂮT�p��x�9�L��@wJ ��d��}�)#n��4�ڃS��=�:�X����r���k����ύ뎁aa�BKo`�~������7d���:eDj=ss�L۲S��BQ��-n�ku㒙��^�s�]�c&�E^W!)S퀽�y�s�5&�'�""w�Ko0��*�$ܑ?���lʴ���mtd���j�Kf��p1���Z}_i�M\Je�w]XX�=�7�J�R��)2I7r��&�;k���H���h�x�'��i~D�[Z�j!����B��F�[� �D�w��e	�'��(�e�jO��6*��+���N��8 Q�&�a��&Ҧ��{ۣ�;��p�u������ԷX�����v������G(�n\�݇��C���k�ϓ��=J�.J�Z��2���d�.bS�b�'����춱��3���k{�v��}ԶY$�$EJc�K7/����N��I�Gu�?���#���R�%
edj�u���㪓��>��ڥmo`���[�ι�B�o����Fq\���T�z�p�t ���Ti�&�7o�u��䄅�9�\[��]���e�ˇ��o��q��nH2�ݎ��܅��f�b��I��C$:�6=!)z�9�s�d��?�܆�W�ܤh%�|����R�Ϳ�.%�R[ØU�����yf�0j������e��j�a�"؋{��}��,膂�` y3���n}m��<����{T�@K�ׯ�5�tb��r��yJ@B^f(1/���B?�Z
�w�V_{r$a׵״ԕ�i�|������a>���Vg�OKN.��G���=%���.>>���J~���ᡴ�Lkk�x0�_AU83�l�O���f���Y]�PXQ��^w~�|@#>^N��#l�����s����3���\L�T+�Hw��z���?���?
�!*���.V����z~d�Sc��9��oOM!�ܬL����vK�P�~Ů�4ZW2�H��jE[ß#虀��ݷ_�T��^H{�l`����k.��_-��"�����|�|y�����<1e�jz`Of�ɮ��,�ͻ	����zv0pߒ6E?��?�P�*���~����~xk����h0�0h ]�s�}��s��ޒ#W�cJ�I���#X��g���R���X�����2Q�
?3�;��pw�#}4&�&3>����sa33���}�"��������Ea2���Uo����l|�Ƃ.��jĊ�@�vG*Ed�os�9�څ�l����d�^p ���g��B���m%o���LZ"�R��u�W~!9�����=����v�Ff�1�So�i7��+�0��6��k����d�W�_*A�i0��O��Nv4羿'm�Ub-\D�Ծ����K�mZy��/ ,�_Td��bj�fxb ��B���^1���Q�h���-XL�%7�)�1��i�������8�l���OOh�\{ ��Sw���ysǀ����Q����gZ^�{��xMT<�<	�-6��'I�;X<��~��\�TY�Mg��Yͨ�J�%�l� �p���$�����)�o������]��D��eK(l���)�&���I���o�L�z}}���	1	��'*�;v��Cܾ��P&�,�9���8�8?}��+U��MF����H��3/�~��f|�&�X�lB@f{�;���;�G�A X��~A����m�).�Źs1:�_c����������ak�ɽ���[�r�\�H�O�}�8�k����ST�a�t�G/]���ĕX�~V�&@g&e��C,�Ȉ�{�Ģ+-Z�|��:W�SW�A?Y�w�J%u����r�G;>��{I�s&8j���jK��&q����ή@��6v�f6f���i|u�mykF�,<(ê�]�4��?�o� ��G�}���gW�Y�I����d.N��:7��:낈�%��`���Q��e%���Tt	.m�z0�Ƃ��ʸ��]旴��G�BJ�I^�����<�޲��mص2-	@?�+��� ���|�{2�|u�>)&
M�`���g�:L}k����-�#�f����k�O�r<�H-��7�Ğ� lU)������TQ
8%�z�x��t�gR���{��}r�4�+KĔ��k�7�$Q�/>�Қ��9W�告����~�UC�	{$��L�%=��ߙ��.��M��Գ���Q����U�@ݙ;:����a���T���B=���n�����.K���[{��nb��Ζ8�� /5�7�8g'��_Zc�L��.#X.6$��XV�Gɽ����?['U�
n:̫.1���q�(q�ynz���Tc�����!���R�ѯ4��	w��:�P�L�:w�(<�U��\!��/�R���P K�G���!an��C�XCJv�I���k���E~e9���B/uǸ��yM?��L�	pq�\Z�aJs�u-C��j�N�1�C��b�M�6K.�Ő�O���Zc�5l�)�T�œ;]��P�D{�y�y5�2w�W�Az��گ��pF/ʜ�X����@����E��u2X~�}ł���h7����IfM��7��<�/G��6$�
E����<y�~��%�׹g�<��/&���#���X�i�!Z�BJ �Ęť��߰�r)�-�뿅t>`Gↁֻ���1^ab�����K�	���|l,���7tŸb�k3؋�F����س4��G���=<�'�OK��ūR��Ox��rP���ǝr�g�{��;<m�k�����ȶg߾"jG29/Қ�I7a�r1b�ݜ����ZN�Ҫ��ޓ��\vm����),��nR�/q@qd��4H�	�f'�z�'F\���TX�q�2oy�����JZA!�
����ի�H���W����/��r�'J+���C��RcH(�u�K[<e!ca��e۞����ãǱFsΗ�-�Ce����q��+��p����5��u��u�8�w��l�����o:d�_�<��y����4�W5p%*3�\�7聍�w/�|�g�άύ��xq}}�����N@'Ͱ- �8zaƓ?�����~Hn,5���!XcY��aW˸H��-���b:15,wŭsE�}|?�),'�*v�w��	K�����Ǖ�l���T$��dq�2�~�VV��ONK_''��uz�X_�*:����a�m!?#�z�q3���5���G��q��k��6�Ć���I1��O��$��G�`Ii�?3P�����_mX��&���F�?�bG{����"u��N��@r��q�!h��������f�r��G,< �=�g��ma�3�a�B�;�J$�z�^������\��=Kr/x���>a ����xo�}��*^��٭'���ڔ(��G2���"����&0}�a�i���x�4�[�3�f���_�7w+�P�>x[S=y�
�7�گ<�!˃�i�n����F��$\0%�&%2����ª܂ZG���g�$��p%��cVI5{ ��+g�1m���#
�O3pYUFXW�Ͼ�=�X��4���{�чxZ�ƒ�hƭzh�I�es�&�l����ݠW���^�N�2J��)Lw�+��K��r������_�]�W�`�;O���-�3U��~4��X��b�M�f���bm��BR�<�[9g�L��r�/˂������MQ���r4�ť����J�}k���o/����õ�vi��?	�� �2C<t��a�j&��~Á��-�d�kݗ!E�<􄆪��d9m������+*�:��V>�����Y�Щ�Tϑ��9hd�7@q-��7Y/��_-�Xr�Z��]:,GFb��b��oS�\r�Vf��v��p�x(��c�r����JC�o��/9Efݻ�������yy��#���7������^o��L�w'�O��"�T���*�G����
�C�'��F��B�b,j�|:�#N]3#�ĵ����=��ψmӯ6��\��X�kt�I�9�~���(5�N7a?{9DuЗ�lX�TY0&��	~��Ux��ֽ7&�0C6�UY��Wܼ��6O[#dd�����	�rZ(_7k�ÝD�;n;���K)��B ��6�[=Eg�h��	��3Ew�o�o�Q$�d�#��v��g���/�����B��̀��z"���d*����5��r�O���Ar��>�h��n�����+znY��[LJ䕺x�*�/��HW�!M+;C��w��y"��@vl9�+�Z�]t���,��:�i�t�T��%hT�ц����<޻t�T0Y
�H�-��\�8�$I/��j�l1K�����'�.�8�8D1>���޳��~>�`hb��;�'�៉w*���Q�30:�#�P���
��p5�Θ�/]0��p�:C`M�����2���v	��ω}����)U��nR�Q�&����T}2Q�ր�X�%�� A����k:O9F�[�d��$�-�u������7x�a�O���l��t���	����E��'��}p>�+�SA�-Q	���:�Q��{���gn[�OD9e�4�@N�-��7����l�r&���݃��q�_�����Nm5���)QzR�z���q��v����%��Ǖkq�Ŗ���u�����Y�Ý���mW;8|�Uk�r?`J/����t�5�!��9�A��=R���jϾ�8�c�ӗ�;s~p:��V�M+;[�����Q�4�5�>�͑�d�ؘ�����BLOW�a�z����r�eѣ�a�����;�B���/�_Ƴ8���|��K�`�a�p+��C5�D�n,9ԋV�����6"E7� �� �|W�e8c��\�F��-�Q��T��&,4ڗ���F�n2׶�w���Dqd��cߺܟ��u�L��90S�w0_׮���e`ް?c>_�2��$��FL�ۺ���I4����a�/���{}UB���$�.\�B�B�vm.4b�nUd7�A�w����In^���p�c�4/#&����LLM�s�*��+m�0VQݡ�b�l�{�y#p�����U&kN���Z.[��+h�&��P�KK �Bհ|��[`�r_�[^>� ��13[\�G�����3�5�qB��������^�x�|���0��z�98�X:�RE�,0b0t�����+;<^ݞ������Q�%mW�A���=�a�+��&ey�T�pL��uj�m�t�]����`F �������ʠ-�_-AE����I���!��ꝫG��k���َ�%p5��9��6��'
��{8��{u�����)�^�TNӰ��Y�݋��:	1�ޚ*9~\��8�8)Ҹԓx*��ah&T20xv��o��l.�ײr�����`od8�����ug~75a5a�~��^5[�#h���Vk�C�p������8M����ұ���`c����z-"��-�)+b��Q��H�	py��A�ok�:6_B�8],>�l�<W���Z�5}��7n�u�(��**�Y�S
�̚��sܗ�G^B�}CVL��&@f:I�Š�#�� �w����Q_��P-�-�D�v>��Bι�h�vx��FZ´v��J���w��9����!q�N1����d�ɖm�6��{l���}������/����^n�Q}�4�����+�M���ye%^|8I��	[��.J˳C5����fdD|Ik���dTdJ�J�E��~c�g�$�rHZ|I=O�@%���ճ��`����d�u={���Õ���k:K���w<7G]��FK�Xx�L�b#w^iLJMH���G,�x�(�/��3���jLC`�Tv�ElAS=K,XA%me�۩w[�ɇ󉊮�/�Y�ŦG��%�yg��@�������vP��ᡗ"�i��Ɩ�f�Y�! �u�Yd;ē� �;�]py��~UN�]�F�n���MM"H$�@�C��|��L��
'�}4��V�������ʯmeQ�7,x$���kYٝ_�J�%,�(yI���|�Da��;�x�G���Y;�$~"�. \��7�#�=��J�'�]㧷���G�ͦ�q7��R�O�n��|j���C�ƣE�dq�\���'�������O.�rum�I���첞��T���"�Ăr��H�$rթ��Y�!����I��V$2
���G��T�YOʸE��w`��h�=X�-��հ��Ų7����ql��0�T(s��q%#���>����[\�M{����>��Q�6��<Ii	p��7&
��[nh\c
[nk�����^!�~��s��J�MN���� �!�&����R���u���	��T�_8=�:^�\����i�a�S�=�MG�N�����ݫ�w����Y�M��<�vO�x���}=�������!�*6*
��g'ڰ�����$�ʶ�sz�}���_��	���(�J�._�ז��~+vCn�z��_�D��Bj�2|+rA]�ƃ�Z�r�N@�>OaG��H����`F�'D�cV��zv\6T��E���t�ms~F�t�=DI9x�ۘ�Y;��1�l�vh���l���D�:�#su�D���,������Z�*�	���X�e�T��l����'����ԑnCp��U�~��WF�_��6ˌ->&�M��/[�,pi*--�U���Ը	L��\lm0=��t(�Դ>L�b�Ӹ��&){�O����6u�>X�SXޔ��������?�S8�tf�S<e��������@�3�ג?)�ѝ��o6	=y����x�'�����ϧk|���'���C"��##;��qSMyyy��1W��6�e�Sl�6�1|׬c.*���:����-�D,�t��> .�����S���'��5̜]���d��x���c�u5���+��Ë��EI��~n&k�X�k/~��Q9�6�3�F���M��T{���ԤGC�]�^Z�r�;~�Rܣ�ǐ���_7�aċ�X�j��S7na�Mvwy�w|�s�>�[�����Ebff�����őL�&)�շ5� ��f�<h	��,&`��Y9��=���x~y��-�y��^F�y!J�:���>(7<r*���H��������d0% ��,�pC���P�F/�f��+��a��z_��&pP��U�qY�I�/��������J����c4�93a~�}�Ō;8���;�p�/z�M�&�uч^�������>����{AsːG)�y��۷m��x*�**.{bZ::�#0����q�rL�] _^�_�6�_��ډ���T����ߊ��qb&��g��W��F2��k�#R�h����?��8�E��y�i^�L6�BlA�y�<�}�K�[�Z�ƨ2�'�pE�Y�^탆�	��y��J�?m��ף�OXG��^�F�6C��ֳzEEA!a ��>�J����9��i��PkO�AрU�UT���(#.#�Zw˙��%G4R��y#G01�"n�b�?h3�Jɰ�v;�ִ��=֍�.3�G������i=�x݋v�=>��ݶRv&�2`��g�}⫧]����F�8�J�u;J��$�.��2=-2)�g9V֩u�3����GI����L�o�\�8�u�I��.����\��m��M���g~w��d�E%d��dڀ)�M%����t> �S�l�������@,#
NdŸ���v<�d*�qQ��M#���-k��Wd\��O&�/���<.Z"RW�����F��� �W][��Wx���e$H'�T
�s����#�v%c�pct���=|��`�����Wƃ}'�y>t����,���n��b�o�ESc�d�|�M�z&�oii�Kw�=a%9�Û"~{(����K���(ْ��]{a�G^�ˌ��ͅGhC-��@��ˌ}Ï�`^��^���H�N�O�>���9�l�qC!��~'����"��;:Q�zW�r�ܼ�#�����E����K#b�`D�'Q�����Vx��Шk�Q�N�������H�;�r��4|�a�#pB�xE+�����o�*�<���_���⋷^�������XT�/�;{���R0��D����\�k�T�E,����s���:�L��YƯv���m�8������ѧ(���$+% ��;�CڹSr?��mo�G􄰲�6?�߭Ơʾea�'|���>��[�q#o�+���no�)R��O�~,� 7�A}���ea������o9���3����MO�����bPt��B����}�3�؉Ա��5ރ�9�$���u�CZ֒���e��q�t�=z���}�UQ��/�8j��G�|^�C������7�^d����I��JN7_P! RT���$����$�L��Ҹo��\)K�������6R�y9yK���֗��4�Y�3Q	ɹy�kV�T�eX�[�?L#!��(��t#��ݍt��t#  -�1RCH���R��!�0�������</x�u1{�����Z�0z����D�	0g��S��xTN/��sO���_���%��_mcJԑ���X�N�a��ٲ��HhX2��I��@�) �)}[�AFۭ��kvf.!���Cf��ٮ\��t���ɗޚ gL��&u��Z�q��,\�����mi�B�>��Ij�H-�(�<�rF�Z��aj[�Tڗ�D�S��;�F<F��I���Gp6a�A)NO~oV�����Z�t��Ѳ��>�vP���;!��)}���Ǡ�A��D�cǏ�;��0���%����WrC�����$��X�xM#P���ޑ��m��0�+Y��g�`M�}���-6���H�B��}A���.�)�.�1µ���$�>Z����%e���%���BA�丂^�T����
"�yo��YܢN�<���rÔ&�O��s��{�fS�}F8� �$-&ZD(���M��蝄j+%�w��N�#���I�l���0>���Z��=�(�_s��~ �d��2�C#��sh��?�T+b��_q���Bl�r�I))6�}7�K&��=AZ:	S|�!�6�" ؝lO����V���Nm*�F��P"�����D�xla�naI���Z_2��D��CJf�}�6�/M2={��h+���P��wgdA�jY��{tV������S�\_�ם$�[_Κ�]LⲆ�����ҫ{����Aǫ���Vm�R�{�%
�n��w�w4�������b��wM�L�h�8�g��"M�8�ӠT�	�*�v߹�UZ�<Cn�uy��wa��B�{���Il��т�q���6��Zoy~)������/:ӊ ��w��X���dX(�}�w>?
�Γ xq�����uH*�P$6�B��tR׹�v�*S_�����I�D�>�����R���3��r%�6Ɲ�@�KS���"������ə���-�k�P#<<>p���ycEVX�#>��pk2ʤ��L~�Qo4^�v��� �����ʬbt���²�`)��N�Cx�kvO�lcy��@�k0	�C��Vt�H=v\���CK=�0v�jJ0���k��+��	ӂ��2ؘ�~�D!�n4#��6��;&!\vĈd�!gp��#V(�h�5��0���Hz��'B3�+r�F_��>9������� ��-Δ�W�����ǅ	��N���������	�p�f[��&�T�;�_~�x��;���3j'�������Lac�U�ͼ�}N �+mϏu͖��A����Rm3�B܄*�Ǎe¹�e�o717?�>�_����c����C
@V�K��|D#S�̌��J���3��`��._�W폞-����nX��D���'���\�n��bͻ�?��5�?�[.*h�t��֖-odK�)�%-�:lJ�6��Ĵ���4�g�薪L�I<��}�B�A��s^�Zk�zE�C���0��/~�p�z�V�*��n�S��¬�J�Q�����Ќ��!�p����ö���5�4�%5~F�.ܧ��ݏ���ܰ/�+����ݜuRSU3hi��B�v���ym!~��Cu�X6���'n����6iPϽg,|�E+�WZy9C��f�<��x�0nQģ[;__��Kf�������&��Ć88��&��`�D�6����5�ܰ���Ү�������h�p+������1`��[ʡ��MwY�SK8�G�xKZ��J���	Ji��oC��Xp܀ ���#�2^�t��V��[3Z|m��NҠ�d�(T �z�;���;d����h����שWֵ	0:U�5��o�����KzLo[N/�5F�`棵����E���Gy��y���E�'&����0/�U�_�	���޿�:T���,a�L┽:-Ҷ�HIK#u�hE��8>Ͻ�@_� ��GT}P@ �2{**��b��'����/����&#�a��6�ؓ�:��tP�ն���U_�x�6N?f%���hXz�bL�\ŷk��bǁ���T�˷��f��������ߛ5�����pt�$�_J;l'_��%E⓾l|w�x�&z}+�;4�s�\ƿ��=ƛ_myR��P����T��?ko9�~
�ǎ�b{S���FE�Ђ�f�JKK�W���`���}]g(��'����A&�{��י�i؀��d����:�1��:V�2��S�Db�d�	��v�[(yg��J
�t-���'���wD���Z2��|":��>�����Qg��6*d[�'�Hg��PS��O�^Ćap��� Y��b�^K�䷟d�Eք������VA��e��G}��O%%��4y����?$�g5��Veى����gi���t>Q�cTQU;�Hb�� ��-'㐤���|*$B�/��<��e���d$RL!E�I=���pe6�wR@ޑ��a�p���[��
}�$��o����5k��@���_��Q�p���0{�*�Q"aH-{-�T�K�=K�#�����%z^uj}��u�����ЖE,���3dqc/)�^�Q�7�;��߉���������.���N:��^�f�G BO;X����]��./�v�h��soP����'�;��lo�d��:��$	qh�y��L�	����?H�o�ۑ6��x��Rc��ǃ���G>=gq	-��{��A����ނ�[jē� �T�ӣ6�����q�J�FX��ף��fU:���?��w�sr$��]��d�B���J9R�?�x�k����`+�������ǌW��`�j�Q��a�Ɣ�Y���[��8J�O�� ކ]��ԢR���7E����~2+�������I�Nr��O~u���O��ێS��IQ�[�E!fs��<�㎊���H3){��&�����L���x��܉��>�	$}�����O�1D�ͨ�IU���zW��{�����2u��]O3��u.I.Þ��+�KPH^͸�q������8�Je�9e�d�����j�[��Z]�ͯzS^��g�F-:���U�X�a����Sfp����
=AYٔ	7COp��W�d,JJ���r�T��8����:�WFc\���sr��oz�MY;?��L���{��u�7��+��L�3�C��G�<����寒򵎣�� ���w�Y������w{�)�GK���R�D� 8_`�c��Q�o[��r)8��M@�3�������»���� t� 7���1�������fB���Q�����@x�0�߳��|.�,hL�`���ME�B�	P��{w���V�j�t�X�j�c6�[�?|��֍\�H9�Vs=�	�	���BM/���큖�;h?`81VaTZW��M����T��.�ݒD(��0�盰�N���X�>R�Ѱ��-�6U3�b�@�*R=e�<���~]���05��wFvw\k��2�5k��V�L$��~@7����j�]�y������Y��������"�66X�&���MV+�u�L�2��k�Q��"�6vv�����@(�e?Q	��񉐭��J���fS2$�eÝU����p�����q��k0���	ц]�����<1E��{n�	��Z��AP�s{� �L=�b���rW�<��~����>/�u�3о;9���3.�:^�d�$��+�9��!*��4�Iԫa#�k<����7��j0��R�:C����7�}�X�FF�$���f���.a0?�Z�W��
Y&��3/���jQ�KR��'�Mq�~1�}Y�`'�OX��Py`������2��/EC���W#������@VG�5y{�j��[<��}4yQ,+�_��L�;˦*���{(7e�hODc�R	���P"�O�!�|+`�7h��o�w�!=���.s�4vǄ�!ò��(��OL��2Ѯ{.a���R}���fy;2ݴ��e��[��l_��b ������D)/�e6�e��zT���آe%���q@Q���I�f�WQ��?ߵǔ���r���$%���9�k��V�d�w !߻�)@�����~���U����m���o���fgz��7��3��Z���"qta�RR��I###t�H����~U����'!)����������{�)>&�᝹:c�FN|2y�3p�z06	����"����B1̒y|��*�H�}���o�X�d���6��Ï˥��Wo�zuT{we���<����d��gJ:Q��'�/�"^�kf�N�v�c�+~���|*����^<l����v���.���m����dz1��Oѳ�'���]V�,�\���U��J��$�W3��5��3E��dOP���x�sV)�Ϥ$0;�yn�(C!�Yp�WN�t��=
*8|u�<픤o� �y�:��Ȩwa_�!^,�׉kp� ������ry�8��%�5�
���\:t�����R)Ļ�~�&�bT�L�V�"��_^h]d袞�Iv�S��B��Z_�2��#�>א01�mX�k���g�=+�<�p,��E;��@��w�����¸�/����I�O����k:�H�!�xZɀ��|�@�\SQ �lmm%db-�������|��\X ���f[�Fyr������#��V?�Lv�@o��������݆��a�{JL�tFz� ��Lg[�'����NN���M/��k��2�b�7t�h����,�E��S6��Z]����<klP�>v{�8`��=��O�E}rp�n�_�S��{�j����J�/B�iUu5؇��p$@�m-���I�)+v�=�X��Z�'�0O2s8���D�K���ۓ�m$�*�����F��O_z�O��\�Q��DI �* "�4H ��qɳy?^���]!C����py�uǽ���%߰^!QɄ��[[�)��ɓ�I�����Z����~5��4G�j3,��t�t�Y��O�F+������㟭k��cSS����a�p[q?��D3����+��Zfe�+�Z�fD�w6�s�`�a�[z<#�:�����
o��G�_�����G��#�Q�a�m�b'����%#�F�1�]*�)����A��'�!����0�����`۹)�����������7�!����]���*\h�U�)A�ɻ/e����l/�׫�����@<?#EUE�9�jaar�yy2�� --X�P�Z__���.�.��Kk����{�臾��x(|A��6�B���e��{���Ĥ���-!���G&��m/�_E���u��;�c`q�LM=�j��	�L����� K�/�n����S�s�ڔ����O��7�*$�j�!d��	�w���aL��'��,����C���O��c	5eN�R��D+��-�3%u��WM�\�8�F:�)z�zwjy1<����U)�U��9�o�����~a�{���y#��y�=�~�'����s��w��d�2V�9Lw���^Q $L-T����]���L�j�vޭ9)��^�P�Y;R^=
���:l���z������I��ex^75���~�Jb���������<0�E��O��{��꥚���ib\������;*�g,��\���ed +X����.�5�r�W������G�6��������/�R�G��~ɮ_�sx����0���d��r�@�6g���0b�h9����c`*�],��0�����3t]��#{w�'Gb����;��-k[eb#�4����\�A���gE�x��%�j��N\�������RM!f��&@��7�<�$pK��b��-�@xM�`V�0���r���崸�R�SO�1���y+o{��)K�����O�%�Nm�+E�3\dW�kΖ�i�=���=�n
��9d��R�i�jJ�r��Na�4��U���"4�#DN��9�#�krr=Fee�#�9NAA�Q��`Gb��L��ш4;<$d��#@�	���b	�}�����e���1�g2�)T�L��HRRk;'��r�Zh�0��<<2���9﫩����㽰;\ � pѦzu7��{m8����w�I0��_Ow6�=ǎ�/�l��F��F2M��p��^�ojf�^����mc�� 	���ڈ��F ��Xr����!��Px�/^�m�;�r�ca ^�� �<a�,���f�m��+ٴ��b�yMW>�xM{��N��HĐ$Y�O+��ɜ5��T���	�.~��S<t�%퍤���}����6_xmooW��3�AX�Ɔ��V�i>[y����v��7<|<Ai����7�4�h���Oϲp��jK��@��u���!;+�/f�/9������=��oE���>��ND!66�c�`pYX�-����.©�T��[@G\�d��S:F���}]����U�%2�5��W�:�`+�w/[ـ_�
'��G2�I�����͕�V�F�%b�Svo�agD$!a�0l����ޗ�L�z�$
��<\�{���!mԩ�F�93��|����T8�V{��C�]/��?۰�T���Q��B�LYYa��+�B�jy����T����M�G�	�#��֝��Zm��p�9�#�>G�wn��a,r�bs�X!#�=>�)�m@��c����%��B�����a� ���>�����)7��3���n�潕�k<�6���]+ߦ��O�Z��55�8�)Ē�l2��P��m7mG7��Z�Q�ЅfGRIIɲ��ψ�'E\D;�,b7��F���u��5fTy�^ASJ[
���]cϢą����5�9 �׭[�ݲE�g�)>dgZO��V�s=s~��_L�T�����w�K��R1=^DMB�1` ա��:SZ���S%%�|ji�z'�ak�U��}}F��el��;�"�D�/SI�~�-�������,���KD�j�}���
�ʕ��5�x���qy�O&�	k �v���g#��ԯvK�0O߻g���x��(Tl�U.O��W��c<{�����ASzG;Q�8�Jdo�}}�=���3��W����>��� T7���f�&`Q�/�]��"���8T�* {�E���Gc�f�z�CO/�>xv��/��8�{�ZUt�Ҍ&{:4:�ibb�>�TY����|Y���6*���-O�p�wm+;;��EC.�����45[UU�< ��yx��%��Dd�\��" l��E˙oqs3��R�M�K�E��pB��qo����s<tr6gz*���=�{����Nm.��W�L
#�Ap�D�1��&�H������㚏�1�gQ�p���Y���W����ܾ�Tl<C5�}�
�ׯ�(ʍ��C}�GU�|v���ztG�]f���i\O0�"���6�`�KLW�Qn�βC�綌sn��M!O,\�JDWk��R�S&��-�7��>hu�=�[�Y��&�ޯt�ȷ��ҺNgf���X1�s[J=[j5/̆� a�0���� ;�Y<X��8��ώ����T��B�;+T�[�`�-â�&6Z�"gqf�>������a�������Y�p��� R"ù+5c����c8�&A.�C8��Y�_��+�<�M�!�����@�p?�d)��.��v���������"N����j"�]�⌊���;;���I��|��ݩ������h���SWG����5`��Ğ:/|���	�;�k��#�3�(_@��B�@�u�����Lx��nq,y?��ο=(��6��iJ4�0�dp�.��Gk��\Ȇ����,ߣ���ӗ�o�L�n�Ok_�/[��4$ y�0�NǃZ�xR�������ӊ�f�.'!�{V������Kl������W�+�3��T�;/�魥X(�s7�yl����������ؖ�ص���,���n�w~2��U�����cXHt���
���Bd]uף� ���p�h�D�_B�V��m3[����OԎ�Q��������X��{�7�r�����i$����=Q������D�Ǜ�+D�f���;�lV�L�
m�D:xV'2�V�W���WC�����{�w���eb�/�������,y�0O��1h�Dʟy�(o��C��M���S����p�0��nQU�!pR�3f�8$?S �Y���_+�nIlf�o��B�"|5c(���_'o�aJ嶚8�N�9ԏ:@>2���(�鷰�8�z�����[m�7}�cr%=��k����Ӣk|II)F]�!d,���w�+�at�M�s�.2��5���VN` <t�pi��soមk[0����߫���ҧ�_�/1Z�����K
�X�����!�@~zs;Y�]Jŝ�#G��������i��C ��TTT����WR�'
���D����k+|&��L��f���M�ϵ�8�ͯ�04�Z�����l�m�x�M�l�/��^fe������;�e�\ާ�;}���z���i��zB���?�O��z O��Wi!�i�}V�c�8V]九-�1�_'i�Lj}CA��!�;� �}]%ů�\�Y�=3��9��n�j����Q]�*�����G�}�F9C��q }���T.AF�'ȃyڃ�p�_�F'���O׮���Y�r-�vҠ|�3z��&,%������J[3�IVN�8��b�ޱHh}��n��dG�u�7�+}h'`&��հ���SA��c�R#������Z�@\�&�g��F�c�[;lv�Uƾ�_ 4(�B�oY&����F�:��ޖ6�ܖ7E�܇:�M=9�ȏ���`�GL���T�9tI)��M.����w&���F���nM�u����x���gAPWbA�e�3_�d[�t\��O�c0�y��ɬ��T���g�j�M���Z�P�������Y������X�`kW����Ŵ=��v�^�9�z���u�l�R�^ژ�����%�U҈��d�#�q���n,��oP��G��ƍ�����j���Eg�n�<aŕ� y����c� `���v,���2����&���{.K�E��q��'F���2��8L> �p'*8LqN���1�*5g_Î���<��}[���
����,��=x��1P�&eb���[y������`{H���ac#L7����'��饈>����.�XTi���Sצg96yz�ƓP���[Խ�>o֯{�`pi_�#
��j�����\ScRXt��6�s�=���$۾�f�8j��SƸľe3�F��Η�S�Ь���"q%�?�@yE��b�B5 4O���IBϥ�Y��刯`����{���U���� �F���t���/l�J�قf�^��s��2�L]��H����/o�t��|-���(L������дq�^��4�U�?J�gy*�μ�}`�W�|5zKmcbc�Ng�ĩ��) {���p�r�i^��:�=��9� ��IJ�ZQ=lԩ�<��>�pʯ1'�b���x1TSF�O�3��)��}�kОM�����R�?��'/t�r��7Ęo���S\�ש ��E{�ԯ~
{�����w�@���G�2��N8X�:X�"���'6vKO~���U�۝�d�^�����)�.�d4�o��/��ܖ��'�^0bE��e�[��fl�!H���7�ӏ�[���z:n5��7M��H�r�vk��;�����{��� 'Veoo�����a�_O%&|�9- ({�;��^�v<*��{�Z�
S=����ݓ)���n,������Y�ۻO|"���AE�WB!ɇ�h��#��w���c�ںl_Ӻ�m�R׶��@?�ig��%G�X��U�pG����ZK���#+?~Q��S.� ���AS q9.dH�����H���ݛ�o���|���@p�,I�{)O�?DN���8�I�ox_8�0�=w7G�eevoM���wM�x7>�W�<�=�Y�������b��'�grl�,2(�3��::����c"��:<�yF�C���o�0]�!ߟ�\��	=���!6G�/�rFq��Oh�Z���a��TG��g9sT���[��9��Ɍ��*�rm�tC&��z�[���a`����	�q�Q�P��)���|�k��{�p�6�tg�z�����+�`>pw}�
�z��gNO�z-A����>��HtTvR-�n�� �j���Ĥ���:���m�ٖH�~��8(���'Se
R��Fz�e(-ZR[$�YP��`T�I%�u3P>Uu�2,��xb�_P$��\���U�A�N}����&�/�>�a�Y	:*��Yy����kۛG���(�¼������۷��JY]�l�9��h�|f��&��Y6�2�wq�8���ĚK�"\&���ߩ�^�������=*�u��N�E]�E�@�����ͽ%>'�FVo|�U�{��o/m<ݲ�_�Ϩl@|�2#��yĊ�v�N��!���:���O�Nt�4���Z�\����wkFB�Н���=�;�t�C���E�C�����������:mtz�Ɖ{���mh'���C�\7��Aq��wؐ�������;5���y�\D�?G�kQ!�޻Ab�6���j, t4U5	�(h���_���	�pHߺ�1����	��Խj�b8r����+z2�GEA�p�H����s�Xs]��}�gR�mPG��m��s�n�B�������ϟ�m���9�op��$.�y����ָ坠L4�Fx�e9X�F�hq�ӈ��vɴL7%�v�/Ci�� �~>�-:t�^d�Q�HS��[ʑݧ������_��B�8��i����Ȍp�黿��^`���N�4�VR��U�#ď���8<�)+�vIe�O}=�q��8,���A��#�#��V`וM�xH+#����A�R��z����y��L�Ċ��]4x�9��ږ���uG�E�ތVg�7��8���$ r�螯?{'��6�|;[�cP.��(��h��/�j�oku��
d�T�}����m�����3���I/M�{Tz��)�?� ��3�Q�-�Ɵ�A2���i�
� z��)����PMOg��&I�a[/��_��g�|[,������p�.6!�Ch���x ���D�`����B��cߧ��'s!O�{[kʩ�:ɞ�=/	\���vJ�����M��}b����z���ug@?�NB�ރi!�ߖ�U���<g���v:���/�m�݌I&�u��充[|��0)�4��(�~LП%Ŏ5��F&?DxG
Lo������].{p���V���WٟxcX�j�ƝTQ��b� �П�X3%�V �3�8�&<Zk�D�,���l�uT�{rd�DY�� {V������2���|N]�k8�u�(*��[#�����zqj�&��a2�y����isr��W���Ϗ)P�1e�U�����g/w�?����LR��(���2d�����C��_2�Q��T0J	w�h¼������~�x�v=24�r��EC{�����w.��{�P��������+�$���Y���ӎgY�:>��ue��¶1՛1�"�^���%\~Ad"�7]#�ȭ(���	1��~ݴ;�
�ZI����5��]E� ��]'6_X�AY�=�|U0��d��:���݀��i5O2��O���[NE�ZY*8׎��/�:��a�
����WЀ������[�z�O�SLI�w�}B����c44vx닐r2/�Z	5�*�^R)~����~�����R�=�G)q���o����{���=*$��_5i"�7�-%goܗ����lr�KN�����Z ȗ����t6M&���) Dǰ�U8ER�-�`�ߠ��񫷟o�m�g�Q�2ӳ���8C@�AA�@
z��H(s�Q�W0Ц��	He�� ű��BU$�Z֚��U@���_<���p{�(���N�ޅ�CKwO3�G*�1W5���A�&E�������)�������kL>�D�,5&��z�{�-6�^�>YC2�w���,�×[eP�mfoǢ�
1Bd��:��?���~L�OKVnؤ�U�E]���܃m+s�0��L�<�����3&�7�i������Ͼ�x^����j�&k]���|��>$h�+y~мS�qp*����T�@�m0:JЇ��2���[��)�kM~���B���yG�M���M#�����B���(٭-�ɋb�e-U?�{%���V��\�.=;��m�����2~�T��~<��L$�g\8���Z^�69L�M��c�B�I�]#��!m#�σ��)3_����vE�lk����q8س��jV{�\ʱ2��+��x�.��������K{�Iar�ĝA��B��1���l�_H�+�ф�곲^=1b�`�c��_������6� ��/X>�V��Uv��-o�x"4����4���&)3n��(d��B�z5�>s�za-�n���&gq?<�yI ���ɳ�#W�H}v��p�V��i�W�_}���99��n������tϭ�I�{�~��t%+{P�u�V/M�t��4��w�������S�ᢹ��b�4,�S��^����n7�鵫�R!��?��M�|���Jm�Rf06���{C�s�4iD��=d�6�|�sص�T|f�Yh�ޒf��K�+ف��|�{�O5ܡ"�?uv.�߼>h7��p�Jr8�Q���<��$����i�7���_��J�E�ռ��c<�	Y��V�H?6��5� 4|�$s��X� U��#W
�)c_t��8I"vū� ��G�XM�쇮Qoh��\k	���;��Q�.���@��.d�2�߯l3���e�����UkM3*F˸����`��wΥ]@����G��;����o�Lw�������v�k�I!�1���;ˊ\�hS��j��<,�R�p�N�e��Ƈ��˖R�0��!��}��Q$��[���Z�y��ҭ�8�r}����0��mʤ�@y�Q�/Q� ���q��c;�)�9>b�gP����މq��
C�l~��d���d�i�6��W�=����m��c���Ο>|f��ܬ����_���7��kDav�)ᵅ���g��BBdzN���h�ke#�7����m�\c����F)��g��WU�(�'��:��+;@4��QK>�[^�d�Ur'�l,�N���mp9iߗ�c!�^lc���E:��D0u��@<eS!j�o�0L� h̀c��_91���	w\��  ��Y�H��z='�ZH��n��|Oh�`nr�yr��^�nHҐ����W��*^A`O�l�Ƕ,�pCyEMQ ���~��5�կ~�Q\��[� <!^��a�y��|y��)�b.�.-��"?���%�e���z��� 5���V;{~*8���
FBW[��S=@�3J'���U�	��}��YZ����0w��l$t�y�q�b�>�B�@��X��+�m��}]T��M)X��K���r���h��|���Q���{��g<�ʝ
�k��A�>7��)QN�V&�ט��>�N���C%%�)sn��wk+|чK|�jٔ��f.�J[�ЎUe0��a�������>n�q"���pws�Py;vwE;<2�-��ϟ�^_�ȩv�F���e�O,�~�������#�ͲX(4*����k�"�@���������f7Ə�K %�G��jumF�/���3��/;s�Hŝ:N����|,�/��E�s���~�?�����ō���L�4l4���L�Vq��t%��P�q��W:`�x[q��.�&~dY��yՔϚ/IL��5��T�x �"}��/^�����.y�%�fZ�s\�Hp %�	�>,��Z�yk���ׅ��2�4ǡ�|�?"({>  +a�=q��H������P��zJCf"�nj[�5;�;?�J(�m��ƫS������?1�#�
�#����`��+��G~��5|!2����x�r��Tɱ��tƍ
\8���lw��R�͢���є���m��DVN
G�;�kg��q�	�s��\/E'�(�q�RΦ=��7Mr~]+G���?J[T%�7n��{��$�3e͐>�k�q����7��b�2����iW�]�(�⠳\�m" ɗ����߹�7Z���F� �+j�(l��c��j��L0Nxt�4�`��o4q�ڦ>�¬�q)l@D@�FqM�zA֚���(�\��eG:�{վ��30��Tx�{_p���wE���X�*(q�kW󽅳cU�r���ٿ�
Mʞ��*��	NF��`������F������dd���n����eP����w�S��߁@GQ��:UW�����������)	�Z���x5%bfG4�5A�!8CeN�~��?�z���υ궊2P��;F՛�7��vN�����<�����L��I[^q��tKATv{���'[�iF�i�,YF���`Sח�ɏv&���rOt�X?��aLa�t]*d�l0Zv�W��A�A�L�L�`��:ڤ(P��~nE�v��1;�&6���J��r"
�`n�T.�u�}�k&Ch>�*�k��e�U;+EqS�Ǐ".B��2?d !BN?�;V����2y���W���U��>���q6�qy�1���<�\�0�n�aLaWgv�q����9�����.}]!����\}r��)ͣ���=��j����R��	�V(=f<�k�fA�n��Ι.�U�D]^C$)$��o��{_MlL�dwJ8h���F�jia�mu�j���Z�2��>����F��^`�9rPӇ]����*�
�1]B�a�������Lj��f�:AI��ON$��6}m�&d��
�u�*s������cb� Qo�t�����R��$�f(��Aa���o�j�+M5�*�oh�U�g6��jk��qZM�?�f�O���M�������'�F�s�Y7͵�8�_����jܶ�V�G���ݡQ@����������h�6���>���6�={�u}2�2�K�U&�����bE��F2�%�.�-W�I�Y��dDK[�֭��1u��r�u��Q��և�||:c��/py䵚�ij��=���+�A���]'	��2��#�krX������e�_���-����u�,!m���(���(�����!R�aYki�kly�'ü}bT�������c��7u�'��D��	�ix%��+�Sk��&� )�f�&�*(&%�F?k^�HD&�Y3B�qtys �e1���|n����®�����o�1��+��;ٗjj�{X�c�⟏0\���)^�T�̗/� ����rW����Q�D�$�n����}���m����D֋��O���k������X6�����(g���<�����l�]?���4��O�X�k˶
��0����E��q������?Ǫ��C^L�엔����FU-H���y��thp�?9�W���.��B�>o�qb��������j@�f�p�]A�� DC�����`���x���ync�z6������y�4��_.ڔ���{6��a�8"Q�L��#��/#��Q�I`
��g/��������<q�I������������^�a7~f/�g<�Pƽh�=��-������T/&����u��z}�C��J��'��?�+���#��o�JT>e������m�R�r�[�}U]MU�i7���U떕d�&S�����C|���~�T�]Џ�?	���)�r�7�4x1��������~QD�yB��i3+�fd)��C�;�	�݀E��,i` �s���{i��7��?[je$<S���cY�`U�׿��*׿��c��9��*{�aV�.!0J�g#�L�V��c:�G�**\��(^o��(�հ�US�J��I� uoE>�	�F� ��f����ui�h���o�q"ZחE�h��ZK�΢+��&�������T�-⫔�1k�K��S������>��78�lvll��'�ITܔ�u���}���TK�fvl�HE@Q5��d	5
o�d����5�kQ�֔�Rq&`)��mT������ݗ��u��w�{��J�q�7R��A����X�7%�� Zz�������2��8o�ɻ�]C}j Ǌߋa�hqF%$$Ե�+<
����i_�wIGU�\�!^ғ�M�
{�~0��uB��඗+����T��a����$L/g�3�a��X��� FھokZ�N�n�K�A���$J�v\�n�l�� ��KGf����{��2=�S6t4���u��Ń6>܈2��t���~�<IBdtt��،ŏ%;$|����a��'#{k�@JW�C���غ��?  � �a�Aʹ�R�1YEPX �����K�6|��A�f�\�G��J�����:<�.@��-^KpY�%oou�]ng�&�����w'v�ݿ�'�U�ї�CA��?�[�/%��.�f��^amc߯�oŋ�ABT����15%_>2	�3��`�h\x������/��;^͓������ZJ=#��\��8NK��`oio�h�F��y�+�8Ō2{��"5Z_�(%������}�d�;H �ʞQj�M�;�4���n�Q_����a7��~��|�3��Ia���\���ݻ��Y~�^��✻��W�UWa�ə#�\�ee {zz�V�n�>����G�)����i6P��	@���T~m�BP���ؾ�u���2+`#n Aw{��;���ш_�$2�W��+��X��!毷V/��uK�*q��jެ��費-���.5Yc�0JF��-{1B�
��=|EIIY�o������@�:Y�U�<�Ƣ�m0�2����CL�Cp�mlR����>௦!<�����y�=+Ǵ�QE���zd�� c���:�=��9_�������G*�H}���q��������L]��͹���l�|���z�k��~\���¯�uݒ>׏�;��S������M��ׅۢj�ޔZ5kojU�Q#j����U�gѢZ��,�v��{� �.�D����}�?�~����9��s�9J=_
��q^q!Gf���*Z�_~��W)�CѺ_�-�&$$+�ᨊ�<��i.��8Ǵ�����xs����E{���G�Ը�{,�Խ6y�T�D�W7d圣KA�/���[Q�@��P!��b�Dv�|��~Eyu5"����ۯP��ײ��~����K���Ŵ����觸$6��½(�5��pu-Wп;0<� ap����ϧ��e�Lbu�v���ͺ���e���v���X�#pBh�zlNWق,����O�|�G8
�G�9����Rc7����X�4���uz��Qg��8L�:��*��N����p��PG껕�3Û?ĎX�i��f�"K?���m�J��cLzx}�t��G���2�q��L�-��7�_�PG�����x���0�~-,Th������\���SSs�{'`w����b��aT��b>J*����0g̕�>�es�zaR��#�t'a3�j��N$i���T�mG��>�l�yZ.�� $��z�*�����s�2A�#˕){�X��9]��͘��d�[OHO������AU\�ԁ�I�e�v�<$����2?�����9G�A���R�:��+-$�^�X��������7t��N�v�./���!gڰG_>��>RF\�}�.Q�u��Ӣ�><�&�����a4��f�����KV�l}�TCBҶ"�la�.(�nڤ��%+�n,�~{
[�=^7a)D��L���%?���;}�s���yHQ{E�D"7.��lc�T劌����=4�E4����ަ��>m�F $�n-P� ��c��!�b���r�������)�g��d��~�������踮gl�Z�"h�iQ'R�Iԭ�Z�
H
�g�	��ҥ������7���_�/E��͊��\Fl1%�O�Uf���gS6I��[CZ��}je9.�S�����J-�P��ƛ.�(:L;��E��J:����*�X��^��x�5���Zb�e`U2�l)���T�봸����c����O���/`�:�z�I��������c=B橨����(����g�Wxڟ�$�/H�gK���ݘ�Urjm�L���#gu
��m_��[?��|��[!hZ=NNi1zq��|X72����"y�*���K|��@\�t��?T1��	�s0ӝ���3��'f/2�}g�ZI��K�2�/C�V�"r���d���#l�d����P홍��Y��lgL	���ψI1t^��z]�^zeQ��,!�j����(�k�a�,V|��˨����Q]
� �N��C���*����S�D�����	���s�Z��}��ɟD)jG������S�&�}qs����y��3�
�.���'�A4h����`�j[�k����±`�E��M$�d.�R�����x��B랉S��Fe|+z�����lڂ:E�`�X �qa��g�&�/;���~"/Y����P��{�w�8��fk��yB^N�z����������u��Ie����^���D�����?��66��L�sb꭭n�c�ЪZ�oEd#8+��oڭ��;(��&H̀�;��O�T��
`Ig�2�#J����H��Z� ܰ��:��%������[��z��L|�#��ϫ�N���%D��{�y��jIF����1����oEzb#�l��:�6q���>\�_��`���ߋLD���nC��uk��0�O��.J|�U)J;#n��:��8Զs
���r'ӑ'�/{To�iڐ|���������!���xGT�秠��)~o�DV[���}W��߈�k���1�����sttD1���E^��3��X��y��X�=Lc{�K	��Cvs����#�輻�3;���j2�>k�����`|h���Y2s����KT��+��ȂuJ�4-�[��$Ҍ\j�r��O]�]d�w���!�XVyZlEf���'\��L=��;�q���.cOg���������Oš���.�-��̜-`�"�b�8b�C���q���C�4�B���8;Z���;��f�烼WG)�+�ߋ��L�o�� �<h�{�Iԅ
����cS'w°t�:�N�tu�@j����xsj^<R����D?��� ���W��Y�c����o�'u��
b:ְ���C����۫ߥ�)̷Ǳ)���ψ<�޼���WYƔG��C|��:/�|���U1��[�������8G�z�����o���F���C �J܍�]�
r����F�����k�>��
���'�*��-�J���\&���<��OM?,�38u�e��]E�z�o<j���q�<cˤ��<{Y�]��y���������
l�<���#z�̼b�.�*�x�p�����,�|rK:���:r��]2�+ɓ���K�|@@������S��X���co��j�9�.s��r�)�-�ފ�12������6�a�>������ǫ�v����^֓���K5KtV�������}�pY��?��	���_��y �w�ܤ��.4��{�Zyؔ��ύ0�+��	�<���jĥ42�X����8e�$��ڕ�n�?�l�-%[���֗��I���g.aN�C�_Z��J�Ը;�b1�x<�O�j�e������(�]~ki���WQRz��[�)`��q$S)k)d��|���!gD�0o<]�dwߒ����f���&иf�ēBpڂ�{d���o��U������"���=@�}	��T���=
�s�a0.�)���Ϭ�E(�CNc	�2�ٵ�}���?���:t�DəC����nm�K�<F���0�Y�$ä4��#W?	;H��T$&Yi�_`���'<k/ŗo
"�_0�x��@��<`Y�e/�7G�B��;�/�̷#F���j.Y2h�������6�W͏���ql�k�3�"ޚ��*�)n=�hf�����mI�}ڷ�I ��~���t��������O���������b>N6�֮Yhz�9��vY��9�"�6���7S�'���b�K��C��Ta��魍��=�q����J��h��A�?�5��X�z�,�BH/�^�qD���q�c������C�^�U��Wm���|]�4PGl �hF8����n耒}�i�Lo���G�=4�6ؘ��I��lnT��oG�d��4�oE|LA��Ӵ���.�i��2��(M���ֺGQ4��Ҡ(�eyRo~5a�?˿���0^��\n�+HJwW��_R�Z9`"2ob/���$y
9,�,2~��OnO�m�X��PY����7��Xg�RR7-�n5|���-��_hp�"Y.������L��IQ	()�?s$
M+iL.�_]@���Z�֬Q��u�>%.��4-]���&:(��T�6��T��xY='�S���OP���{�7�ǥ��vV����j8���97t/�hyς*��8��5�m�h�����E4��d���c��h�ѹV|*����G
�w!�$�͗�Õ�{���YX�Vp��&�
�pe-�PDs0p������O6cIp D�R.�(dN��i� ����J�����*S�����!-��䬸1�x�f$��@�mP�<j����%`%(e3}so���������d��<^[�S�N�q�(�:�`N�E�� /�T���/Q#�Fd��G��vա�_K!��T}i�bџ���������ة�y'�
�~r����d5�%��e��F|z^&u����Y����@�ި������YKk�i�6?͙q�x�]�/^S�`��0[
L�/�����* SS�¡�����%^՛6�\F����͗�1�CÂ�(ɦ������%���O�\0�v�A�R�����ӿtc�S1U��P�o���&�r��(PF��*>i�շ��!ۘO���+
�9��ח����
:$�mM�̡���_&��-$`R�f��k]7j_�\�5Ñ1�g������R��[	�gۥ�q	V��ϡYq�!H�9؟P%��2y�Y���~ȺY��OW�vX�xBG��|-T�tY�;���G�l�q��O$�թ��l���Ӝ�l��C{���'�ԢeK�9���f�
x��OAa��Ѝ���)�/X ���4�?H�eJ�r��������� b�#�9��A�[mW>w+1E��u��;��g^�
�q�\��{9����������|���M�' ƛ̈́�u��񞰣Q�^Y���c�b)�Dě�p��E�9ju�GsE�=�B�S~��Wى\�l������m�Հ�HG�In��,!k�f�b�#�v�cӒ}�� m��ju {Vw]z�/qu�NN��&����ZE��O�?���� v��-�k�mC|Y����[�G儙�e
m�f�+��� ��X�N�$������I^A�ӊ76JJX���'�������~�`��G|+�DC�8n��8����Ֆܦ�,N��秒��M�Mw�(�������=�3��-��g{���{��ʞ��bhʤFj�y����r4��obAhf���/��ux]��(�����<Js�]}�2�WQ2r���`#�a�HK���-�^�Z\dpԽS��k�?1�
2ϫ���lu���a���v	6#�C�{���3w֚�Tª�}�j��4�.E5�u��y^� ~FjlĎh�L��n�ΞI" ��,�^�ǥ�]n��d-6�F�~�$����xX�=�^e�dI![4k�3�&(#���πIv�8�Q��:�)->��T�-�Z�h�d{ZFq��T�M����J���je--"��Kk�OB%l����u�N��`�s�$��YKy���Jz��j�R�S�WU���TQ�)��9�S�ߊ��H�3�����f�P��IS~����"	��h��@�o�|�u�_کljj�h)`=�Y�w�}���^��|
 	�^�|G�ȍ}�݌��m�z��]>�D$�����\�СN�ͪ����'_�q�?y�vE䓁DV�6���K��vYHk�ݗl�"'��+	���hgE<%H�F��p�a��}/���ɷY��7��-���������V�����e�����w�{����������M/��?z���j�{;���¯K���&ce����[����s���)�+T��G5�� ռ/<�8���u�T�a�U���g��5=�zWQ��s��Z�9�XH���΃�z�\	�=�\q#��it�^��=a�H��_H�j�1���n�s��(�2��O���B��i3���iT$n��G��л�hʟ8Dl�l�sq/���.���t�U!}ι/.�M�|���2��L�R1���6$b]��vN��Aǅ��S|�4�� ���
�� �=���H���v���[���b̕���1����~^Q���N> p��F6!�x���җ�:�L�r��ԟGȽ�ԩ�R3�� �`��8 �0�nz��;��6@�Z)��NR�m;QNf��~,�ޖ��ھ�dY_x��B���sDD=��W�5�t��D`�u=��I���;_�E	�,���ܚHk�8���ӗ�/�4Z�ih���齌'G�.��PH-.���M~���]hl*z�_s�]kR����O�ݞ�>�L�#�I�k&�-+#b
�}�����Cٔp�5eZ?k����5�׆{��[C{���i-�ʶ���as׷���V����kYJBε(��g�J�DFPo  G/=<jꙋ[��=a�.!���H���;E+��=�WKL��٣����Bo���Vu"��nq)�4t,)L�#Q]W(��ks�8��Ӹ���z���i�2��&�4 �e�E"@�ϝ^T��y�#7���D�<;���ˮ�Q�`;���K�`3l�^��<��̉Y^�s�w���A��k��%_�=�a +��o��%<��Wh/���LE�����
>�o�xE{4�t'h��1/��Z����R!���LY�
<��_4&����2{O�y���x���+��Wl���G[�d����kA����$�]UX�+�%���^��H&��D_��E�Ć9��2�E��qHcu�]��xT�"hY�i���s�ՀvL�It����f`jʟ�r��5|�uN.[�����.!0���Gy�ܡ+вE���A�����;,�!�^�7e�b
yI0em�]5����qU���E/��Iy�R�t|�{̣A��pW8Q~tt� 3�{+!�T�0Ǚ-ݯ	W^�G���<�0\A1_���/��1��})��eNqFb��9���jo��
���p���#:oKO-}���>��76�-8G��͹� ������w�$�
by��L�]݆��g<M����A��o�4E�)S�q�&2bx9	�y����w���0&0�3`X�r�u���H�V L������U�֔�9��)$�6��qSKKIL ¯���C�ʵꯛ������� �@^Ycy^��9��F���Nq}@�_�ܹ,�	ڽ�x�����K}�r��;���qdFF�Ѽ�����( �*�aYZ�$�|�G���%��j����#��'�(�<�O������yq���N*�%hմ�[`�n�番���|�y����G��¡�ЕX�omr��������OH�=WH��v�d������aA��aQ<l�Op�N^zn����n<1����2�?.���|�!�C��N�gi.�m�XF2O�
���+��Z�xA/H��s��҇������v��Q�^��=�5���r�g;c�*���o�	���X����~+���P���C0�-x�@"�籶�͟WD�	^hu0�^w�kV�M*!0c@k� Z���������S�(�q9>�UͿg�Q��O�M��(��cm���.�wy������F5?��`���|�f� �,<�� 6՚:�=�'�2hn��'B��[9�$tRy�NW!��t���8�:�|B����` �^,Qߐ�;����ѣ�F����3��]��ʡ��C��D��c䈙�[�톿u��xA�#ALK�;��Ñu:�à\�Q�N�����j��U�P�g��a��;crON�d��K,+^�,���p�b����.n�z
f��I��E�y����a�U;8!�N�H�o9�����X��ёF�w1��Å^c�Pe�Cg��G���R�^�����n`�L{��!3Z��P����K��lT?HU��^Z-�Z�E(���wg�Y��@Ҝf+�����A���0OBQ�
`RI��2G�����n<��R��G[Ӵ��6��>�c���
3���R)�%�
��C��J݇�R�3����'o\S����0�-?:fw{�q�ס6s�ς[A�,~�K�����NN�!鎓7�L=p�4�"Z�j�A&�˟A�/���fW1�4�v�O��]�d�<���ݧ���xm:���9��^o~�X����*l����,K��v�z�`4������H�j_��`��\����#���m��Z����r����@�,[�PD�S������G�O�/�.+�䀤{��@�j�^�iW�N��n�MY�UN�Eƣ��'����|�m;9�A�c���q��d�ۆ������^mx�V���4b��'��O/��O<�������x��<�n>�]t�L���<�Z��G��-��j���S��_m�x����W�^��E�t<�'���ł4Bz�z�-Ɗ���~Pы��}�P�!1sO��-h����վ�WA����wz�xk9ˋ5����-��
��=���2#�r:�H� ��C�SȎΘ]w��c�$�T�����-����2b�#�O�_I�d�Ҡ,�O0Ζ��;/סLb�ō~���~Do7��x�R�ٸ4	�ͩ�0	И�!k/xD�Rb{��Ίm 3U�E>۶H5�Gm~����9@i��G���� u�͋�� �����侂
�_ BA��ohƜ��.�9P�v���B���a!���h��E4-w<	6�����F�V/�r:�?{x�Z>�a�t4��Bs�c�%e�*ww}����y�*>�C���YsJ��?�\9�5��"���ʺ���姀�]���7T��w���?�s��`2���U���V7Hhf��<�VΘ�:�����!�n:��^��n�Np��9c.���Ϸ1 �2�X0�7�7�Ь�XJ�}�Q�Y5�χ��[�T�jܥ����U����_�ks��k�?C��pDGWF�5�T�*���[�!eF�0T��{����� L�����ހHDkd��u�s���s�o�PbQ%C�2�}��O�����/��,.XHc�+��������_�p�z����70rR>�W��I��p��p�/�C�3ه�)2Qv�f~�9�ɭ��#���83�2�
��3~��D/N�*s��e
�����a�/h��@T���mg���wڄ%X߹������(@��L��`�5B�z�%	���KG�E�|�$q[F,vZFCdF&H����l߅ �;7=�l�\/T ��PЎQ	�{m��@JV�w��"G�p�ۮ��]Z��j|�W��ъ'��m (��]�G;H��2����D$hj�>����Eܗ=����+�/L<f�ct��T�D�GlW�ѕA����ס���Ն��!��E�&_lKF�u|G��8j�|˖X�Zt��&yGE�Q�G���yB�n���l�@�nބ��O�[v�hP+�E��)�I�D���a�g譂G�=S�xE�}�&�H3��J%�O��*���]��\k�Y�o��6np&͟@�\?*L�&�)8���E�RG����a�2X�>/(��2:�	)��|G>o3;	z���8�KlvF?�A�T�k���/���jI܏�]���x��p�׼Z3����U��<�M|#�~�mV�.��	{`�쮊�iӇh!K9�����y�X���%�Ϛ��+�1g�5!%2�,S��s�Kd�_c_��>OHK�:6����`v����|�h�F�e}�����}�횙88�"q����zw���Gd����g��	!�p�"��w��"��@k�(��p�m�=::�=j�'"�^�M<M��\\�����&i�"v�K�̌g�`x6��l���*+2+ƾ�͘ʵ����l���^W[݈/#+z^��dN*�/�1.�M����?(����l��DD�i9��I��j~r��.D���!n�#�N>�����P�o�nTC�n��1�k���WPU�OI�z��x�F����U/�c��/��	<ÍT��ւN`��{���2�=_�������^���<(G缈s\.wN�zw����L/5�i��5:����V/dΙ(�ƈXo?�1q�o�=;�����6��=���j��������r[',���-�c��'w��9��_05
m4�'�D�է��6��6v�U:�!���K��Пջ
*[��q,�3��0��*D�q~����V�QU`� ��\z5sD�0i���t�ș��������M��uj<d�Z�d���]rL>>�:j���0��(V�/,��ܥJ�yc#BM*�MA�#'��+�;0�6���[��l$`u1Jdz��2���d'��T����3��~�3�9Ӻ�޲M{��;y������:�C��%����6y0US�H}P��9S����m�����������L��c�贛���n�r��~�j���u7d_(�Τuq8R�c�[J7�#����+0���S�K�ĒtG��@7��K;k��Θ�Kjxc2�sQ�^=^3��q �4���e�-�>����/{�<��H��<�؊��q<Czg�H��9�2?��m�E#�R)�V=qN����T�4#���|�m�M���2�׳f��u�Xr�ַ�F��Q�Ƥٺ%�?^N���[�鄓�^��"�w��^���{R��P�mi?b���"f��+W,TR�M�-Iyko��#8�q�ܓ�{X,�g2�cE�O��ԥ�����hl�,$���*8l�[����~�B+��h�����ᖖh�#�Ass��Åjd9Z���\�VyTN����Ok$�ǎ�?��hd@��6�c%��%�K��cKS4g��M���_��x�AM�������y%%U
o��~yw����'בy���p�jF�����-b����毗=1��%ԟ��4�k����sJg�X��i������ͷ��@\���e�����Eh{(��/�X�9%�#a�a��i5Aɗ{.�M[���U����4���gB�O>[	�t���\�
�4��r ԑb}ހd��o�2����g�Ś�u1��ؗ��$B̜WI��.��
�u�2�<��E�tw�������XonX���Pe��a?vB��k��2����\��ꡃѪ]���<-�6]�8e߿�-ʺ	6&N�[��q
ۃS�b 鋅~K��bޢ�=�> �ݵ�Z���~JD�KjjAG��{��6�|�d�i�*p{���g��
h�E�_�a頬�/�2�(vl��������߾��X�:�W�r���ү�^k)���H(��bu��k��5je�Z�\e�zsX�,e�O�nѣz�}dݼ����4�1|��t�ǩ��~B�&u|���/��_��J��,��~W�6�՘�M	*TP�W��Hw~��%T�FDw�#gt�� =F�כ*�>��2�l�_o�F� ���~��ʏX���w�I�����SA�
���u\�����}��hB���˶�sh/�	������kF,CpT���9���xB��� e��X-��r3�go*z�nN�Kq�)�ѧ�}� �?Oܳ�Nu�`d����u��J?��!�eaz=VnPQ0(������i7?@�!���%noJ�܌��e�yk(:��`\���9�d���r��-�����i�.eޘ���	THS��qx�kX�����2�im$�LƦLý!��ݙ
hm4�G�r�X�>��TJ�k�.�l^���D������Q�2W����nN1�wj��ё�]�>2-^1|�l��W���$Z��6RP�8戮��Y�
��2���Zǉ_�I��8�b�s�|�yj�~.�	<wH�SڱϞxd_�9we�A�9@�9�$찑�ʤ ~uA�:��V�����.[��Ꞔ������Q�4u���gXt��`�uE�|�v�sy�>��l��NNaBT9훾Xf]j�h���dߛ�J�%W�LoYq�QL��6����M��V��7��O/܇�R�9�6�B��#�)`ErL~B�ґ^8rێ:�̿e�5���Gͤ��u�h�*.�6
y�V_t�P�TG��Y73w�����hM5���2|H��$�Q��W 56���t��ڀ�jȔ�,RY�J_q�����1�즿�����l�ighZ��H139�`�����ԈVQ'SYq�h��5Nn����k���e��Aj��ҳ���)�����p���[Z_��p:��Sų�a?�w�@!xѯ�~x@�xA'vw[��f}�Z�W��6�2��=��5*����TIpn/��_8I���ZI��LiPJ[y-�����x��|W��\���\�H|�KD�9��yc�+g�t�� J��Zv�V؆qW��y����-�{N��5���B����N�{Y����a��>��=�����l�^�R�� WS�����Z��a'�"Y�U�����Un"G����5V(\��0*"��{h���[�^�ֳ`ꜫ��'S�/PCy)<W�9�O��
��p���!z �8<�A.�q%>�D	2U�H�{_/ �������1��uU|7�H���W������][CD��������_X�~ӽ(���VL���hڹo;��t��%bs��ْɚ/��{�8��?�y�׷��2=�`��r����, ���M�'R姹�;����O*�2�K�5�����T����bSM����o#��[5����3qɌΉ��j�-�-�9��ֹ9P�Ef�BMҧ5�����hfJ�?&�p��ï0j@_�&�=�˺z�\	�U�����i�b���)=͍��<�a����ӆ�&fyw��<�������:�j[�8��%
�W�aJi�}�]W"S�/�#I{�1�w
���H��i�#X�36(Q��5�g��;��MS��S�.��[�i��^�17>�*�W�q�pz��'���2����O�J��򴴟��9���߯��W��1Rp�_~�e��Y�/����b�/UUq�<V[r��~�J�]|�A�7�����r��s��x��w W2v�N�OZ�������"H�#c��9^����'ph{��`�u�2pk��s����v��*[L�|h����C?��S�.��
���Jf�L����L�w����1��_�\e�t���Y�XU&�pkA�O��;))8��)(i�LBg>ǟ��*v(CE�Ӈ�P%��i�F��⁁�v0Bvyy��� V(/"@���v6����q��;"3�J椗�F>,�M�SغQ�c��3�dӈ��a��9��x�}!�0�镣��C�"9%/L�n@�+�!Z�s�È�Ǿĭ4n�}R�c���Q��ĥ���ޗp�R���Αډ��J����X�P�N
��B������m��<�>��:ZZDttt2}ԟ��nz�2��Ne�|��'Wn$�%�勑%'ߋȫvg��,c�'�!�n:�,^���X����r�)�I(,q����b꩏ÞT���������[_)"�":ucߣP��E����B�دǐ�6G��ˇ��N-�l�*�I�E8;;OJ�S��8����������y�?�����)�Y02�P�]�
�����u���1B^��m��}��k�NWz.E�:j�~m��@^>+s[uS�oii���D�z��p�̈V��r��VY������w6��i-:F.�"���@ծ04��!�@e�W��%������*��6��M����3�?���~�z��rC�|�<zws˖.���N�]�}$���X�sCt@�n�@�y��� �����ku���_��]q@�E����!Q��6�k��s¤|�B�*y����~^�R�'�/OmΘK���
u��*�z�I��J��r���F#���>K�|8�b�/�����f�����C>~�dSW�8�ع���N������5�9�:j�_L�l6��RB����k,������[�x͚ۏ��`��9\'ؿ�jT@���ԴM�D�rʄ����^��mM�\�VL�w˖:�59s�'�C,���U\��7�?������ZX��\(��{b�DYT	�^�6��5�=���Xu,���%�ԉ�2)(������ɥ��*�i\4df���'��<<�(4$y,E	O��Ж�@�7A����z>���M��ү�*ӷ�aG31o��z����� �u>P�gh�0A)?�P��<:�'.���'��˻_�vf�� MG?`r�%�ٲ�ܔ�ebL���I�rJz����!�g�_$}M�s$� S�:�u>3��ψ	���<�qo���+�5m��4�{c$,��861��|���)򠸵�g���p����C���Tܾ"��1Q�J��B݋���R�+��װ��C<?�_C� 3���%���է�:�v��I��ݻ��0&���R)_����@�I~3�pN�r��2�n��Q����VR�#B,2�������WZ:M`���g�+j�NtT���p�3??����ۿ�Y�Ͳ�S������(�Rso�h�2��}��x���\��B�%���~�o8ѿ�s�F�o�o0p�8��DP�K�;'ocJ��lҶD�p#à1ݱ����s����5��\tt0a2�hȄ�8��y���eT2�,����A�P.�C8�I&J����j9:j�{�@g[8�����Wg�a��֛@-"gg��.�T��H��a��s�h����,+�,w=i��>��v����� �`�w��{aCn�|�>��!X$��j�R�^_�e~inn>�f?�0�=�Z1���$�[ɸh[6
��jP��@�����S4��):^,��5������T�[�(8f�:&�4:o��ɜ�G�������8��l���������\�j������󆝰�A�L�?U'bu�!�>��H���)-�7J^mo�S�0�n;��8����F������׏�������3���S@�����HS����b���2�r'�V���69�����ʯ����խ��4��,�lI��0�q;����e��,#��v��z�ؚ���U=���VH�1��>�JBӨ�E9"�1���O�1uj��ɛ�^��ĉn:� `v�|di���(|�������'_�o͔� �T�|e�@{�LY)oI=����B͹NN�u���ޒ�������4��w<���������������2�@�I�+!T�������C�w���=���ze�h2#�X��,�F�݅�-���Q�.��D��H�ׯ7��m���7�/��eS�L�,����]��/(��� �|�|�E���+�w�J��������v������P�<���_�]�~�/��s��5��x�7m:i�P�P��\Z~s`�#`��F�N6��c9<�nn0�%�ܑ?�{ak��Q{��_�*:�9���m�X4$e̚�H5��fHf��g�ΘŲ`�U�-�.`�!�v�ɓ�Ց=�����������޵���AB��E������������_�ޟll���)jhh,,����bL�b�X�:����8�u���@�^�e>�-sj_�g�.��cR��:���Z_?��,i|Y:{��?�������6��6~�`P�7W'j��hGZ��
�����;ao����B�_bW�����������v+���������k�p�,fo&��aї9�����%. ?����c[�-m��Fc�;��_�[މ��X;�R�����"�R�~���K���������}mov��v`s�@�J��9��oo��.����9��ʜ�>�"u�B���+�J6!u�+�w+����W�Sȷp>�<�JP��x
[��;�jK���Z���2(���}�$V��S���)��f~��^�n����ɸ���3�=��bQ�^��>�qb�� �bjF۫P D�k�6��kZ�<
ٕ.D�5cvC=�����d�/"�}Y�����[Qɔ8͆88�r�XI���U|&�2�1,�RP�����
�>��i>�#E.��؀���z�ʧM�U�~.��K;)RJ���1����b�ڏ,���qνec\�c���n���P3&�1�Ҝ���\�2�j�%pJb_�u�{M@�ʔ*�������4Y=�<�?��4���y	b��5�������H�<�p�|H�s�|��v��D�wvt��� �j�ϴ�f�� ?�_ҲI`��U,q����﬌R�UN����?�o�s�|"T�C�i�\Y�w	��V�81�n&Bٔ2��5�6��	R��9��Ÿ@����`��G��5��ŵ1`#�d��h�K{Z�fA����V�Dr`ܙ��c�T����OJc����a4�Xm�fƽ�r9��y�*>́+����g�&�g�uǳ���#+i&&YǃqcUs�@��S�\�"U�s���7���&[r�o���@� � p�2�/�ӛZ��������h��/�"��վ�M�ٍ�@�r0y|D�۽r[2Lv-rQP��#G.YQ�������ߺ� "�s���o5c6��~�"A�O��Ȧ�qQ�������tqU�_SJg���PsF]C��I>�k=�2L�D��0��K�'�b+3׃�\�nT������P��-n�7�b����E"[�(2�Rc�K/w�?K���c8L��@�����}4�8�e����3Hz}�+�֭!�� ��Ds�����©;z;��SĠ(f�`�]+WlƎ��H��G0�
T;Rm�hr� �g薉d����0����K0�蘧�$J�:�@4o�bnC��?K0U�FoV���M��@����~�9#M�?��̄Eβ����'|l��M����	w�9����{� ̰���OJN�����$1]�THg�)U
�?7�6p;W6�F����`�+b�g�r�ǭ-aeUȏ����KWg�!Xh*�fy+�&���|���{3ڹ�zΥ�*B6����4*ս���k��'����	�˅��/�BeN�fҿ�ɣ�3�4H�D�Y�| u����$M� �������wk��]����$G`g�����0�(F��Px��p���@n�>TaÖ3�P/��ɡ�d�^���6�����_ƕ�_y���G�3��� r�C��,|ϛ��w	��b8YI�Z
$"Q��'^7�X�s��Cy�	.�,��)ۭ�m�Y�$ޤ���'�(��]v��=��\��?�x�h���b�osSKwR�[z��$�������������Q]��sZ�^�E&�<��=c3E���ʟ�&��~��o+�ZZ�39�[�6r
�tDD�>���oֵvE:�y+bf5����}^}�a������/7g9�ƕA��n|O�|90����r3ʈ"��ϝ�CP�՘��q�3��w�y�F�՗�x9M?��v�6H�O��N���Z^�Ϙ0��*+%�Z�`*��K���P<�C�:�7.�;��lĤ�Y�Om��1�O���ED0�N{=�m,��u��k�7�ρ;��__���
p�#!�t�����Q#�2㖘�C��"{����_���JO�u{�9x�ɤ�a�����W ��5����Cp�Cp������ݗ���K�]���	�o7��^=��������眾�}�)���<-V���C�p�R�0��`3����g@��g�,"��/�H8�����$�J������(���He�Y�nv�"\�8e��,{e�5d{����7�I���
4�n��@�����Z���w�sҺ���_�؄���I�һa��I���5�l@:������?�6����I6�߄O�����.R���7��fbS~-�f`C���do����k%t�DR�0y�f�r���@\H}�N�KB|�rv`n3N.)��gf�q�˰S"�;��?�.Z���#��r?gB��:�.��_���w~�*!Ŗ+^r���l4B�{��0�Q�Bݞ�Ľ��m����gƯ��b��w�|̇3W�Rm�9n�lW>�F�!*�w�&~��}�ڨX����f� ���h�q��?T`�LOǇ�e<[����o7�LW.�����������nñ�*lL�Ӳ�˽��Ł�/	�p6��p`��z&�7����y��k	�E� �A�<�FƟ$�Hї ��(��+��B��B{�!�ş�33A�ӵN/���)���%Z9 � �5���iݘ����R��kU��I!��Uӳ 27-Y�����5��KO���ޚ��\�UV���׋�#�3����J<��3w��Y�+2p�#��%Pr�5�چ!��vKO|�8��֧�6l�;�ZlF�Tr���fI�	[�B&g��!^FW{��d��罐R\s@噬C��뗆Dga�:I)�,j��)	��;'������rw~��+d��g:�(�1�����7l�|?���jo����cc�ǹ/�J����r=�w5�%�N�DW�nȺ�������PY�7(7SGkʡ�l�c���K	a;�!�`S1hw��m�*c�0ºI�J:\i�u$g�x�E�Z� �r2�#^]HwUgQ|:���!e�Z�p�3��q`Rc
�3pV���)^X�рb����f��?f
z���ڎ�5��w��*����8q��u���m��Ib$�niiD; p�]՗���|t� Ff[-ߖ�lX��4����?���CY['���>:��ӵa�@Q�_.�35y���B���g�L�(log���oJ��{�w̨w�$*��ʐ�n�PW4)IV�f�V����_'w[�����m,��V�>�p�l����D���J:R���W���7�B<$v�/b;�>���~���Х}��W���o#���5j�/��N��Q�2\�`Zx�����r �'Ț��AN)4> S۰����YfYa��MRc��t�ZbTV�S�}�h}�a(�e�~ȡ���)����ř?�CU��!a�8��H�,�]��2�֨�����qa�9���K2�D�m�:�t/R3ݛe����"��:m`����
��_-�g���Y$�����Α��bv��R7;>uc��� �7@����U\k�>��ў8���Z�;ߴIh�r�%���A������-?L���;j,/,�V�E�'��ӕܨ2=~��h'+��g�Nl�?l��>�7�ܱ��W�P�DCC��;B�<��r�����4��hDJ���>1_~�5hM�]k`-H�m�΁�	��VS��cI(���	�� ��I�f��W^���)��G�_J���g�ڽy|������� t�z"I���{�����p�����I��t%D+���ҡ����O�}�7�o8���A#iK�6�C���*�\��&���吖����Ď$�����OeC�O���|au��sc�\)�a,OGL����m4_W	9�,�ޥQ����Bj�r}��e�"Q��;(��o-���|+��Z�c�����%��O��YX�Z|?97X�t�a�}�>1u���R�xk~�4�ޔ��)t`�Y}JCy���X4#�k���i��_�Y��0R��e�״�4��Z�!J$/���6�L+��n�:�o6 VB��!�(J�P�Ł��)ѿ�:��ąg�`���Q�"�0��G+Ni�h�zl�S�!�%Ov���5,��ŊC��P*��uo��]�<���!�Ǘ8�V�����6#��]]K����c ���Ku�^�'��ٙ�n������^�R�ꏇ���3�%��E�tv�B�Yr>��Q�Br��
x�`��9ܪd=��JTdHj�/��c�������v��t�P��ׁ�u�۱���!o��eN��--5��V�[zMw��QS����K�w,���I�O�IO��_�W1XN�K��t�^�U�Ώֽ���*�]������L����b#c�����v�fyb��ٟ�2�:�4���f����X�=Z�������@
�,������(#�]��c�^`�zR��`����7���QL8�U\PŷN��!n���O*��Y�>�}H��z�I*��=< �����-?k��$��x�/����]���O���s6�J���L?E���8��
���? ����wƺ�cO�5��gLNB0��,(���	�ׯJ9H'�i�w��0�#�>.�#�%Hn�n����|Oօ����#��啿�/�����~�k�X�>����z�����h�<:r5��ǩ����~�h���+N��+��ǘ�!�qcI�:܉䤏�a�4	����V�4c���C�;�G����y�!���X��y��{g��<���|k�U����A���,����ȞVD��s#��A~�,������>�j/�\��Y���2��OtG�ዧ&�>Gse�{Y�NGe?��e���@	�����Uu���i�LF��v�9.�B +sVY�lR䉅N9����h�!�G?�7H�P�=L8:Y>�^-�ZW�,v��е�8S�I����깛��[�����'Bt���Fi4��כ�U92���f���Rdu�7@!Ô\ta�?�q��G��w8��<9I8ć�ꑰ�l?:IB
�=��΂QX��0�����N)t�����j����27R�-͛0�I�c��;�M����,���s�#y#�R�.�C��&��r����&������c�?]����mѽ&twE)Z�"�(�g�9mCT4P`^��h�5�/����ZM�Z��-��E?'Ӥ�^��%��dt�M��N(�|i�q&=�i�$V�fd8����_��:]�ȉ�},!��hf0Q�	�|/��S�w�ǡ%m� �@	���qxtr�ޝs�J �+Bvu�rc�*����q��[c���6$��EMY���@0�����0����/w[j�y!j�|d�r�2∌�Ƅ��F"K�DQ��_��+S����V�pF\A`��	���D���ջI�T������<`s�ͷ3�B$��w�:*#��O[҉/>�ŪYf)`֏�j�\�T~�1QQ�G�����f��o/�W��+
�p>��[��m�<k����x�L� ���)��␠�^e��C�V�u?��\�k�D��t�pe+�\�����*y0�W�c��3�������"���i�d�R�~�������+�1!ŗ�grY�K�:�BU�Q�Ws��2��G4c�N~S�L5��[��($���+��N��Q��R���m ��x��f/s�;�O\<���h���n����#��� ?���eտ�`�JPs��ԗ�tp~X?�ܰ��,c0��K0��!�� zˀK]��+JĎW�|�b�ss�2o 2ڧ/C^�](.]��Ѭ޹ɢ��ӂW���u�0=��l[��Og��wv^�8���`�Qv�؟���\`��UCzP�Ҍ��r���r�#�k��H3���9����2E��'~k�@W%�SLS�}ZᦑV"`��6ZS�u!��ߠ��*�f=�������~'�
�A�@)�k�F�}��k�{���؋f�}�H^~v��U$�ѺN��D#[A5��5�Q3��C��q��wgt�v��o9u��>��=-E�/Hg9�u���.�bش�fE.�K�!��ŀ|8-b�7�X�9�j}�˖�������"���*�EG�؅�������2L���ˆ���߆"U?�%�����ᬥ4�Q��/��rPR�qq1-�W��I�y��TxY�p�����6⚧#���l�k?��T|�nk����P`�]D�2u{���Y8D�d+a�i&k���F3D��T��'����	��.w���FB0gJ���j�
��2��.��*E��G�\��(o4�*U�z^o�>�Q�����
����O��K��6}�ڳ��9�Dl� �2��󅩹U���0½�4�Vces�5NgY����T�Z�ttML51%\�Q�nRe�KXbᛤD��x�s��'��q7G�,���t��3�ճ� ɋ�=��PB̩Z��Ω]��=՝|��ԭ��T�������Iq���!4ԙ��2d�0c�-'H�w_�M��Kc�wsh��cZA�E3(
�J�)�0J�h}����5�`#8ӑ�M��"�^�|����t�x�ǋ}��b��Qk_?������055�}��}���=��^)��y~�1�jYQ��U�P�r{����KKu:]%>���n"S��ݤ�HN�-|����1ٟB�����ܵ	��gXHG���i�|�<4
�~��u��iA�o׿�2�#���ޞDy)��t���Y��!���62D��?l��o��)�� �Ռl�ܔ�Z9!s �qZY܉�V�|��eL�u���EIw�v���姵�m���� �F�-���X`�ky��+��]UK�_��/} ����o��/��8�gEo�'�vP8��sGt�!�?�I٭^�?>!w�co�ih\v�.������9�����$��#��f�Њ�0 ��%�1'a+�*��]��"��W
����IyM]�I	9���c^�y����EE�J���������33"������~��@R,�,�۝��`��U�jD懗�h֘��9�v(�Ҽ}#?
Ӽ��#�7Uţۥq���z1�5��ֶ|��o@�	���X�ZZF���I�Y�Ʈa3ӈ�غ��o�#� �����J���n|K�O���?m/�X�����y�|��s?�x���;�aҌ8��d�S�ݭ>��Jt���,F8%p�
��=ɟK�aխ�Z����jT��`�n��r�pn��/�κG�΋���qޅ�г���3eBV,��ֻ� ѺWɝ������0c���3�����ď3|���鯛�v�W���Ъ���GCN<X���k��{q�##�4;������}�e9@T-SGI��;��?�V�Q�|���|��og�G �Q����ew���~�=/���X�hx�o�O�lT��N��ۅB��`fј�0��Pղ�Y�=�Z����^9C��t�LߙZA+
k+Ԥ��`�yY�B��[��-.<+`��D>l�e��N�<Rl7ٴ$7�<[�"�O���t�Djc)`$/�'���4I!�%,>~]�Ce;���6�QU���(X��(7��T�\!N`�U_~Q��������3c��W9��!��6���*fI�4�7�>��n��X�����>.�:|��)��������.��W���.n�w�z�|\���`�i
�|ҫ�dA�����0t	^$���_N��l�d����@^ir<�װS�E�(��4�4��9�w����s�_��:(��b"
b6/�_uUF�^\z�珮���[���A��]b	gH�.4}po��ܪ���n�}�k��m������0�5�����s"�:=�N1�6,�Ҿ�`�v�g4�y��yl�N����_!�,�s
���3͖��S�	X�۳�����5�����ι�uo��[���ƥ�՜[�Nn2��.����EV��_��C9�Ɨ��H�D�Z�LL�'o�d��nd��O�_p�w��bS�r��}R�4�7FE�e�{��Sb��ik��6�\k�.��*oC�������
�&�g��������.���N"6�G߃��jy��qk
-��fw�?(��P�� 0(�u5�k��iw�,��D�꯰Q��5<e��I,�Y��6��<z�@�A�LUM-��j{�đņ��൘e�Q^�</��\2�a-E�a_
u�&��0�B_ߏ�@x	*���3ysSy,	#RM����/�`���BKl��+\�t��
��{1�&5[$�z��ye�l�:]���2�vp$�Q�O��0�}��'��б���6Gǽ���~���ʇ����qM�o>P��F-!p�Y�W�H��`�n��'����ΐ�1���6����A0�~�H�I!N�uҨ����
�YQ�򡘜V++���UV�k��շ
�&+����� ��$�[������&��(X���U���Eu��B�IL�O�d���j�PC\XQ�j�I9|��&�l�*L��Z���n��ZN�j������
�rՖ+iH���w�6Y�a��ly�ȹr��A�8*����]���E��h:��K�H$����u��Ch���(-�]��R������D�N:��*QN��s)Rݻ���%�l(x�ߟ)��wvB��A?c�2d�do��u�::��qs�0����Ǭ�~����&�Ƅ�3�n���[0�^�:�_�IN�X/aw���y�#���Wn����f�S.�Jެ�'5�������\f���wG�'��y��q�X��oOM���Q�����,�����N=pE�Br�~�n
]b>b8�i����s~糷G�'o��b��o���^��Ja�&Y�=�k]^̾�{�@�("'��˭z"ڭ��ߚH�Ρ��ɥ�sQV�i�����q'��}�$��[���ף���TD���c�z���}p7�Y4 {BԜ��o�v��~���g�����VJ��W%��jߠg\e�Mx��)�����"�RA��< m���@J�f�A��h ��W�ZXV��(�"|F��F��B�H�9r-AD��
꓁A� �����R�>�vb ��b�(j-=����޴���}yFp��N��d��s��M[%v�ַ72DjPbON��)k�DT����,E�H��=�8^�t���?�R��� eQ.��/�eN��N"f�����2��+���E1��#���'�H轤ω,�*uJ��Y�*b��p��vu�3���Y��Gfꉽw���n�0�[#�8'vs�����}�ý�H�` ��m
l�:�S�W�.o�	ѷg"c^��4�H�D�T�d��ѕ��$��ͷ$��H;�A��������M8�4zH�K��g�m��1 _�u�{�)y$ǜP��q(k�5����l#�V����y����H�́1����V�����@��@�|�&��m�w� �����6�;��m2[0���B�5@nln&~�Ɣt!=:�-�`M�H5��16���ףF�2����]#�hƑ�iu����588���XJ�WN�w�gνʉe{���E���@ �9
�&�\MC	����PCn��r��J�j�B��j���zL�����[�(Ur���)3Wp��R���u;>Q&c(U�(�w�.F"(�{
��.SSTt�9��������^�e��P�O��Ӹs������ޞI<��#B���QZH*�j����$�
8�,öe#L�R�9�%KKP��	|?rJ̈� '�ٮxgN~��p�]�X|O\e�ǹ�p}�j�W�}���:T�QZ�%��uQ�}�(��!-Qq{/����eMǰ&�z�-]�e������8�X�ˌ�|��`�<��(�jf���^$i��#!�����Ʀ7��^�ˮ)���e�:��bBPwwt�	��7�Qv����*0��"0n�&#(L����N1]CbL����bTV�}�f�I0�}�R�0�3܊�P~�EG%��R�:x$UT�G+��ܞ�ɪ%�l�i'X���U+�,�21�Ƒw�ߖ�T�X��L��3��%I���aq�"Վ��UR������͐>:��:�t1��~���k<l�&��.h.0h��,i~��#��N�4�Ir�ΖZy�671J��A6j����H���n�4���և��}���Yjp0t�^:�i�K��&��L㧬��i���Ox̪Rh�Q �.�.|6(> W�p��hG���=C��#����@mx�5'I��>ё���9�a����ݟz���q����Y@$��p����چԣ$5��1�z�z�}#n>��i�@UC&W�RQJ`� ��#�E8�����&!���	��������	�.Q�qr
�z�{�������L7�}�?�ǂ�@@�9X
�����s�h��JgՏV��X�����M�'�#�'�9{��ju֚C�!I,,[�{s2P������Ć�U�X�̉��+���
���Oϕ/wRP�����Q�_��*8S�BS�U��b���P86��� w���$��'Ȍ{�c7����⪨XQHu��7�o����C,������J8�ǔ��?���VG5ے����0�LM���}D�?#R[k�A�'�-ނ��E�����G��72ӥQ�̇�?���Jl
cj�i�ƨ��m=����8�q��@'�[���~v��	6��n����C��p���$�ؔ��|���ӣ�����] -��ڊĞ;ؖ��l���.�HtCҸ<R�4Wa=4@*_P��Fm�Q��v&��SK�I$�zg�P^�n"����m��r <�h�"v���/�`KwBũ�ՌTfw-��wҊ)�~�߼��W+���$�+cq��ޑ|������;~����g�{��}]3۬�#h�'��w��s{���)�����8 #�R�
�t�WW��vQ9�x�¤)`��$v�mL8�{g�$![��{� X墲)�QTS�9�~��צ�`����T�lgDϏ���AF�0��
ط���k��c6�{���`�����������/���.|9J�4�r���Fb�I�Me�%:���0����r#�])��������F�{V�����âGӭ�5�V��;hk9Y��hnۦ��E��!�g�,��>�o�2��Fʯ�G�>k�:�t��Nnմ�L�[P�]��3ɸ���a�p��߮Tօ�$�q� ճh?��+i8ڟ(����$PL��G�_{�^�i2~���(��G��Hw1��S��ف�M��6�G$T����b��#$ 0�n>�+͒Z�c�:aݺߚZ�+�{�(D�u��|U��YF$HO��TEQGR�.kE*�+n�f
ڟ�t�;]��h���,ڡG!�3�\�.����dn���;�<�֫	�:�'��}q��߼<a	�Ka AQq}5|�&ܰ)M��H��DݻS[A� �:���Y塕&�/���̀�o�������?�Z#�W�ۍ���|�����eO���?�$r�M:m���"R[;I���0Y�\�B'��$9Am"Q�m�'h",fԥLA�:��D�δ
e�/��� ٌ���.g;�T�q%W�OU'�O}�8��.�c�yn�����/�13y6B��CU�Xi5��#m ^�@� ��㶄����O(����J|�iWL�c�ۦ������������p����w��Nz���1�K�����E=��}jJ�ǳI+�f�P=F��ix{j�n��
��*��~V�KFІ���Z��뿺�c 7����^"(y�0�r}g�UGz`�����Nvu%�x.��a�����p{���6�>8:2>�~����8n԰��ķ�����g�5��! p���������v��Sk�z�/_AӦ�(znQ�� ��t,؄Mx�ݧV]��p��K����p�_��qҍUT�7��Fj��0XF7 lߓo]��r(�3Y_ޝ¹�n�l�(�o��چ��]�@�2Z���({rf`�2ع�[^|�'����O�וE�a7�c�K��k���@NzX�6Y��9_Z��!ߛ�:�ڙ��W�hy�$Í�y<�5������Q,������k�H��}I����DD��b������k�u�'_%$�S��P-!�G�] �WJ��~I�c�/���1=T�C���8�J�s�dℭԞҠ�v,W��<����Ϫ��e�����w���:��ᄢM�˗����s�rKI��C��Q����'	C�C�s[Z��AUϡp�Sx�S��Vh���!�.�:΃��:���-�8+�o����#�Je|�P���dl��ZH��m��� 3/�0�����m͏��y`�G�`�iz�!�KA����P�����<��"qC
��q�تP�6�'�8O.6+�t����]S��UI��XX�Γ�ڛLd.,'
j�j���E�R�t|���xN��kB7Fq������MQJ���dI�Cgc����~��k����o[5���AA��sZ�u��)���O�9�$J��P���A;��1��Tp��B&���0ݳݤ4��"�k��2�+(�&�2��Pc=�����A�	�wn������F�U��O���.YƳi��#�r(��/j�o/��r�6Y}6�Iμ�	�n����a�U�Sл��B��╨�&:�`�	 ��<kF�?ooo� (��d�J�<�lo`B�6���󆤽����g��"4<>ٰ���7���B�ͯ�v_�[-�F�|��u11s�Y�6N���B_�ⲇ������Kl&v��ˏO��F�/+0#����a�/��M��]�.6πgK1�`f�+������t��0f?�)��W���Ĝ��~+T���}k�ة��8�jB�`��2���9�N�Є<d��z�s��}�Q~+:u�5J�d���5�����-��r/�ۅJ1�\�[��0�*{>�_�M�������5�=|�i����~1���af�Br�(kX��̍��E��oѦO 8��Å���P�����Bm��(�������X�1�����������b�Ht��9�iE�\���:|�T6L-7R��_��^�,ry ��*��Y�����b���u�Щ4`n+���6j|�t5�ͦ>�6;���bz����������{m��Q&��H�z�7
8��bed������u��ԁ��l¥Kܥ^Tҷ�5�����(���	bB%�$�
�,j�3�z%v��Ln��:@���??�б��ڡ
�yP��)�ev{REG�T��a�]l`�`4�7�PzƋ�#��ԏ:�~h���df��w��~��S=	x��#�g�"ؘȖuH(#�c�P�q/�����@��3�	�c3� �q���gX|���%�6kZ�����Q��0������&	�����<dt�}t���y}�~ˆe�uy�Y�C�8]
�SΤ���_R���w8v�?!�(^�]Z5S�8V$�������[��q����!�@��Awjv9�(񕏦>R\r�P%��\�[8�mA��I*��У��K�A^_��+3�^����W���|쭟-��&x����z>��)�ŀ2�@���v!0 N����5�������C�[��J�Ou�:�o���H5���X8�Y2�'��]�L��~�{����j�Q�T)	�7����:�jXQe�K���YF�����m�+�kV�z~���tQ"2o��?�M5w��Z�.���~̞�{�H����ݎ^p�	�͇�>�$z߃���f�̓������<�@)s�/ vv�����B��8V]7������Vԯ<��D%�CA���%���X1�9�c(�՘����e�o��eLI�AnV �oʫ;4�G�.�?�Mn;�9�*�R��#�=何=<#�"�?>qpSȰ˫�j��(� &lr橡v#^�RW�]�����b�����Vح�Q��� 9d�A�����R���)6`m����Z��%kب��,
T	š��LT�(�KaCp�|�Ҵw�)t��;1�J:U�8�0<�S�R_��J�aD��o���q���:��U���)��#�4�Л#�E����E�x.��,%8u�S��7K��|�N�6fS��u\}�Ex��K�2h�ҳ��<܍%�=v�p���lli<W��u�p�
[h�"���+-a�;[%�������G�:�8
�~�n2R݋���T�Aq6�=���ȃ�?�I�|��믏�	�Y�:��%��!�fk����c�?�֐&�cf�-�5�-U%��1�d�iF�����fW�k��(�������\Y<���N(/g�[������'��W��; ����ּX����v��W��o%���<�yo��]g�V����R�Po��att��M;8 ��qEW��>h؆���r�����2m3w���C�zg9k�$U��.��6�R�f�`���~1c�E9ǌ��F��V��qKt�#j��iK�N&��Al�h��(��,��Bʝ'��^@��#�B�&&�o�?��W��jQ;D-]���8 ��N�iZԢ�w���Q�`�Fq�^Ծ����]<��3�S�����r
l�(����4f�i)��&+w���@��
2&5 m����)Rp�k+Lc|��(q�O���-B0�$����F��D�p��~^E	������x��|z��(�$db����r�F��AL�Zh������`E�v�`��.l�=*�ָ�ᐠcg�c�4��z�E4#/y�[��e��1�0cӲ}oH
�'g������N$a�p7Ζc.!�P0y��D:nѷ�SI�*j��-�G���n���|SbZ�iV�8a��P����9�CS��*rH]�~N'�>e��Nc���)�$� �`A��05��w��3�*+a�@�+̣e9�Tޓ����ͷ��8|Z�pc� ���6~�W�(�0����U碩Gg��[�875�G�c���d�8�d4��{�>���܀N�\z��a%dd�Z���~���U��$���M�_@�u�~9So]oS��7�xXS�9�8�+��~���&���zp�w����Q�TK�����Y"HN����jI=��0�e�$�P�5��U�⽙�d숾R3`'�.k��~ �����d�b�����隍-���)	{R1S��D�x��^�%&�vf3���QBN�mHD��f�HB�߲�f����b�~�1^ �abbG��@x��l��r8xAB'
k+�?{�jR��<4�R�]�zR�i������0r��F�r�ǡL�f2h.�c�A�e{HF���o�F�ϥ�=7�q�g`���H#X�hG~��0D0qC(�f_x���Cu�H����-��*D�w�D`�ٰ&���,$�@d)�7m�j�5�l�kE�4f?������Jx���{?��Sw�y{����G��s/:��2�FDA�
U�9O�}�ĩQed�~"60n���IB��cq�'o��i	SR�S���'C~������/��� '"��� O��}�CIP�Ƃg}������p�5�=ݝ:���ה��%$�H	H�=��>+�����鉌<�i���A'8�0xi��A*TT��H�g�gl��i٩������D����}�ȯ2�o��{A��+Z$0K��� <�N`����;�hӷ�K�i�Q%�)�X�v?�O�D����6�k�	�����#��w��js�
�����ӆ���a��;#=��8u�r�Ʀ��7���ɸ��5	�%�X)�	ײ��`Z��;q�RI@j�.Z����,�����y��t��}E�����|"�u(��39�>.�����&��0�X~�IX��:^����\E���E���_nnn�
rK��h��Y7�&�3f�c�����DLcV.��!�`�h6�>��h�4����?���\���v�����Y�.(hv��3	Y�0�)M,g��L�_�Z3��B��8��Uܷ<�3�+(�3^^��������:�}%�~#�n� �K|�a�gэ�@I:�T��vgSֳ���t�D����w=J���R�'X\1v��l����_�u�Ng��Cʮ�̏��}z��;(���o���7�vҶZ�� ��9���h�S�z���/p���	�gfʯvZ �f
��뻦&������=�ôQ�·��-킟y�	-N���'��}�1_����z�/��}�_�'�w0�Z��b86GGF������0��n�d���4�?��4k����k=�;XY���������8bm��0l":�ݭ���X�)�ל��-��22];�z7Fw3I�������PͬϨ
����B��G�Ui�ǩ��Y��	��F�%�K��0>�M�Z�`/�?ru���y�����Z�z����N?�f�.r��܅!J�-�5�{�Xx�[��,�G36"�|��	~~�/��6��_�xx?��W##��sarS�������$D�����2�-�]6k"P(#�f�m��[�����0�=0��{���$����R�t��&&�>���։�H ���bu���i{?ʫ�Ӥ����l�3:ZI9鵠;�z�C4����~���Qs��.�&���@��Q�l�H.�yHC��%��& D/���	��P�?���:9 ����\Y�+˜6}oɡ�j�hZ@5	���m����J�# �{��?��wJ��%2,��#(��"\.��?�>��!��]�Gт2�f
M4���%q�H£�1qˤv�U,�&d�oiP�B���Z�Y���㛀�� �����>���tY��Of��q���>55���b�� 0�P|Yh|>�@?��\�j#R�_�L�7k��W>�J�8޴R+�w����+�{xNi�xB�JaL/>|�Io5��H2vz)U����MO�P�/6�7?g�Z��� �p��p�j���)V!	Rd fFp��?����w�����2v9�mD��D`EgǚP�^|�`''�+�\�N�x�٤���~H��n�C�*���q|_sy����VFFO���v������ب%.�rFLө莽]P`z��+��M:�Ɋ�˱�P���٬������]m����6���YN,nU*X�x�ؽ��]+�(�C΀���/��~��̂�k�ݣ1���cvn��!�FQ�e���`P]��C����5A�䈓�OӦ��(���(֧VcJ�>�
��nm�esA�Q�͍rt�ŵ��	�{ew�ljW�s�<��E�G��O������EyF27���j�v�b����
���	�EL���z^_��0vG3�������~�)Dk�T*�i1FF|�K����`�01��3�Z-��4�$4�3��x���W,�l�� �V����a�g�'g;RhE�5V���뫒 y�&������*���J�g��W�y=*����X(��Oo��G���X{a!J�ƹ�F������-0�Pnl�]p�9G�r�qc���&Q�[�������p�/vHG��@ο:��zN;`s\�R$��`f&(������U��	G�|������A�����sk�dH�T�Yѳ��h����l�B'R��͖�im`2��`_\'��ʊ1��˭䀱�fŠY�>l�����ߔ���F�����(�˔1������S�#H��ͤ*T�Ȼ ����d�j~N�����S ZkX�!?'t� �[U14Lh�]413�������7z��B�X�;����X?7�����&��z��Bm.2�Wr�[�.ΒV���zz��>�@W*�G��w��g"6M�r�a�i� �e�����7e��L�Bn��D���ʩֱ|��P��:q%���щ�N1�T���q���E�)~9/��o5�pm�p�Ϟ@�%���"N�+��8�a_��^���~u���Ѻ�S.kE�x��経� �h��Q�[W���U��ce$���m#*}��ߗ����`�-��%�"m��[s=���!<�b�[�OY9�E�R�!� ,s��  bH܀��!2�1��g�������jx��a��5r�1D_5��S���j��ìL\\܍x���m������әx�7��>_����][54����gE�o�7I�5�ꉢ�Z� /k
�a=Ůڰ$?J�{�(]��&� Hz���t�Ő��*ä�KC?�'B�����(b�DjL��'��!"iS��Ϥ�'*��3�2��X�U�@�Pbc�%t�u�)�Kw#�`N���IM�ZX]���˫|y�8��9[Qx�Ho�<\���P�sڐ�1C���������f���Q��Kp��� =�/r�v�A��,�Sڑ�!w�������|Y3v�f[ږ
��rX�\�h-�S8ևs�rD:9 ;����([]����hl3��̡�����nM�p�x�zo�v>����j#�R�W]�)m9��Db��	�sN��蕚��Q<�0.&6�GN�Ȳ�Ϥ�����Y*�
fh��DkcK�y	GG6�]�999�2�1X����G�~��L��+��Zt�������щ ���I.GGG� �f�7bC�t���*D�xޤ��L���/*���dѴ���<=���BCa"8|�ӂJ��YHt����5��x���O�e>w����lcp����)b�Fp�DKf�~D|db�4P�쓍�?7��4A���P�B&�~�#a�^�q�,@��䢊�f8 \`nn���ڽ��@ӎ�U;Y�E��6׫�b���h��%�hj��Gg0��__�X9-�Z�����kT8=_����I<�j��n[�a�����>E����lQ2��h���lV��H�=���Ÿ�]	\F�p0���G��=\;�Tت^T Y����r���ݯ���&�1@�K�����}���#��]�6��&|3�]4��2q�l�k`�FE���s�yH�&\��,��:�hli�l���m��!�-���ڮa��-!��Hw�� ��t#���ҍ�]��i��Mw~��z��C��Pֹ��sE���5�F�33��R�^�&�!�ٜ���o]��*B����I���V�B�u)��d^A%z���f���Jk�D��ν�SY��B�Td�r k��쎑Q�bx*��2��`��Z��v��8��_��BY�Թ���Z�p�2_K�=���{����G���d�o+��\����a*HK��zg˾VYLѴ�nD��3�
���'��=9����oo�oDJ��y�ϳ��}Lҳ���s�YAMB��[W���4l��ݶ�(�0?����W��%f�W �"''��X�����`<4d�勥ا�Թ@��Wʋ�s�����	ּmq��Q���*�G���ŶE9�[�{0�V���_�E!�y�YD�R�A���*�J;��m��rm^)5���H��ތXd*���]}Z�ԑ�9�/}ߗ��a==33���p��Mt6�Xaަ��6��?3�U6� ����$�-Sհ�*��KE����'撴�#N!Kb�gL��j����M���0�đ�m�ȋ��Ig���#W�@��nP�'��A��q�ۙSd�;݀Á5y�X��R�f����~���|I����=��$C���_9qJ����hMԼ���d�Ywi���84$�x��'6��I~{��"M���)��d3RR�ْF���%�����Ȗr���@���a�g�?�LP^|�%����K2�����K*#ww���Q���xm���U��p��p$;��Sp�z?|c�K�|_�^�d}}Q�Y��F��2���nw���R�Pa���a�/�K"ڽ'�]�5[_����>���uCT%[F�F�ݿ���f���3�i�|���F�����&?ur(HduY���2-��X&���(,����'�C'���Hl���O��W��I�-���(E=<��AUm\BWxF+,5\��b�
�[��)�FL����uk�͇�����9Q�2������5�s5��5�:5&��'�ĒVlT9��l�/p6\0��ب�Ă���(j-�1�-��c`��Ы��y�V��;&O`���[Q�r6��M�NQh�������*���@]����j�)�J�J\�����fx�_-(�Ωm���:p��[��Nn֮��e�^ł��;�}E���]�ll5�pr�`Mm�Q�Ɲ4K����vO�Q��a��=����Op��}tq�\��%R�?4-�2��f�7�*�����b[!zhhG%�7\�8�62ߓ���L����q��:OA�����ֱ֮2�v��훹�P��(��r`�}	5�7���<I��BC�l���9�Ρ
�e��zS�E{H�\^K�Ͳ+٣��!3��aһ{Y �s��QQW���mK���9*֨���)Tb��0�{���!NsɆG�T�?��Y���$êx�-N�
��À�NHKcH�j+VN?R=�o���B�Z���ұ�鸿�\~6{#vP�o��4B�#~�+ڽ�/�ʔ�T�?-��*#����{��?b/����+%����Mvӌc`Sly�Dh���xr~>��p�gY4VvX�l������A����D��"�O����������s����
CKY�|":4�N)k5���aq�ט�v�0�R���i�_�p��z{(����°������T*��h�C���:�ۿ-Ҹ�9�x]�ǂ�1�,��_�w�{�:(�Jٯ���W1�TC��AE�܉��l��!VA���0��yo�����SR<k�����P}��d�o/!��u�H +=��r�5�Hݤj���V�|c�j��dD=Z��{��^�����K��G���S�~f馾,#LG��G�|CCJZ�1�"]�G����h=�W�����(����?�����Wl�����Y��q��8����%���$4u&��eml�>��^z��G��|��$W},���:}���ձ�9�zODA���>R��'��x��&�a�� y�0���-��}W�+�p��x��Y
�Yq�ڙ�	k��8�2{s�'�T�P;/�����ϖ<����7bF���5�Ι�fPU�wQ�g-��0���1$�u�gR(�-v���F���{sYD��U��6�hʓ�Uu9!��6lE�䲚 7�H�O�2�����[x�k�jDP����'f�������r�
�mw`�y5C�:�9�R��'K����L���
c=�\��R�O��n��N���^�&z�����7J�t�Г`�A�"�dq)|�o�Y�\M��Yt	XM�A����1ٜi��Q'otDvw�P��ʈ_Ζu#�y�.l�A���?t��!-�	d����"����KP*����w)�㜬��0�����``@�Z���5��_҅���S��Ư��ğ�\LX��H����+HR�b��
	�yA=V�XAH��pz���'������h���2�C �������L[���$*�Ac��B�Tє��J����ug4�l�(v}���y�D����1�T{����{�)��W+�����(����v�o�9j�ϖ;�����ch�`T\���.����Q�y��e~$'eP�Z���瞺�����w�bY�Q:S���
\�v%�T�sRW��g�^��GO�
 �3��Ⱦ�/��^��{dU4�#���g�z�ՈL|"qB[�7�^u�'17x�ј�dC�(]���c�cX���Th�R^���nF�v�rN)��6�q�����͝���Y�$|ߒ*o�`L����>���
X�~����j�5�	u��i�N���HY]p8�I9��?.��®�AA����k��H�P1��
��Ȁ���m˛����o��!�����h��)��tI�Ĳ"��E�6x����W��0�����G��EF����Ʌ�����s��%RQ�)!vW�&���:��-R��I�K*\�)��b�leM���sz�B�f(��,/�ײ� &�z���]��b����n؁/�l����մ|0��ڴϚ;�j�C��:����:���|�
#5�nh�������gZ�E��bU��$,��%�q4�+��F�/^�Ew ��|�B��4���uW��(�ę�ۧ��u���F�3dK|���oc7�/[$]�w���Fg�w!�v(D/�'�o�嵇��(۪+	[��$-CD�W��4]X>Y�h"v*♓;|uV�<�%��-�,�W�iJvv�5�)*��V��7�Q��'"� e) ӱn���tt���t(��ө� rc�Yϥ�����1�D7�ĉz k��v0�w{89�d������2����	+�$%�co��w1��WW,|=�����#�a�kL	
�Z�͉��@�._"xd{e�y��G߾)2�|��􇨼��Ak�c�gA~Hg0�nXs3?PjGBBB��%ةz������p�f�K������a������E>�z���\���Ѥ3�������G�)���3{nͥk��Hz{��TipDD���èV�o�l�x�`�&�M:�e�F6�u����)��Ed7��0����\#9E�X̔L�Gm�)Z]�N��3n=<*���m�1^|�U>�I��f�G�0��V�����~�}gTI6ߩ���}��ۚ��\61��<�=|=�H�0r�I��p5�2�6#FD�k���R�'͍ĵ��ROBBH������g��P��T��{?������%�GW��G�@�%/����8~�'�'ˣ0^��C����~����D���*��I��1q2��(ގ`�:��r���|i�LD��쫃���n͉V=GA>ը]~T�p�͖�dȸ47�E���� ��2�2�!8����!q������Kt�J�Ԁ�mKo�Y�*��|�O+E�`9W��yҊ@o����\䊍	���?2TeO�ДU��b��I�<���Qu�r�`
�]w��i�$��g���F|���ϔ��>E���WF���	��~�DQΤWXlPN�5
Y�A`�N�������Sa�� d��!��kj|�=n��ӻ1�|>l*�t;��H�9�1�pg#�4�r��'���ZHb�ecTmЭ�-�����M�,Z��ap\E���>�$K�~+Y��ѫ��'>(�񉶥�������I��r��L�.���$m��+��{��cΠ��ǝ6�J�����}��F�������v�N#�wz��/*%"���Y��1XIOOҬK�X��`�C�ݧ2�i4���:!���[n����h�	�؃ϒW�N��r�M�B�0ޣ�]%չ��p�`�|����8q<c�/[�P�_��ưP��~��7�u�A�#���q߃&ei�^�%?�@i��FN���������F8-�!uXS��<o_�#�>�]�cQ�E�r��������aHL�~���>_�
<������ W/��pԨ�h˴y� i�lon������꾫�Vv%�IҸR9i>�bF��G,�eפ����XE�S�������MJM[��6��%�����ֵ�X���>&sO���������3wJ������Z
����K����O��0�/TG��	Жؕ�R�D!�1+?M� M�QP}-�����,{���;<�f6�1�|Ԣ�2��C5���s���ۓ��÷�K�Bi�(*wͼ>2�_�����&8p�ս���ۨ��r��~�) svv�Ȫv뱔S㨫��΅6~�=l1�C��2��cͩ��`�vr����4��I[�Nx%���=@m�df�T�nhP��u�]��g�@z9ɵC�Rbe\��w�>�ٶ�?C)�m>X:H<�o�5c��ÌW�����ۂ��c�7���F����Gd	{�:� ��qy`x\�Ƈ�����yf�l��}s�x�{�lڥ}�}�}su�Q��KE��;�����+��������Du���f4�B�ѣ)��_M:ϩSK�2��F6s����p�dd۠Ў!��v���o�7~�H@��Gr�^�O/k��W�%L�~s��ߞ���WE�;��}_��ƴ �[W����+0�:K%4B�X6^�f�{�����#Ô	6nV%�W|}@�o�;Ψe��/#/�a���l�VE5����\���j�i��3OG�;���\6��S���j.2��u�_�/�����w��@�i�n�*Wc;��S�B��[E�X�����vwBlvw)��#&�Q�%��l���{��3{~��;�vE��۟УRNm��l��t���τ�~6,�~]c�{yA�5���؝�3���}3�՝���>����d��|�G�-
�! ��']sܪ�&��@!Ш*+��V�8����e��7vk�A�+$��F��&�H��<�mݠ�hE�W'��P	�n��ݻ˔�}UX�"�t����8�E�-���B5�M����O���g�@O_N�(P6��C�CyʥDX�y�^���
���v��!"u ����9��MOOM߷7�/7?P��G27f�F �p��Up@�sj��b���FB�h��.kEhܹ���dx;�t7<�4�����w6˞��Q��{.��Ĉ19����|\�:��E&��DL����>�=�S�p9�X3�+���8�1�ڍ���<ߞ�	~C��+D��֗�pz�$���x����ߎz�[��ټ�A:k�� pg{#��(o��6�E�CPUd��,�i`�u
zS*W��4v��_���˂���MT�&gf�ّ��X�9�3j�d�>�ܝ��l����%��	�Gy���x�6xG���혁O�q�u�ȫ[84�	�rrJ:q��Q��x@f��d�����	�$Wn����%ڎ)����S�^'�n��L��-+���:�)3�idE�!)˺n}Xn�4cM��4��di���)�	����.��� �-�ק��lv���^)�ڰ�_��$ �/�)]ۚ���VP ՐׅT�}���n0~ty5?�a�F�vye)��A&�o����N0Eq?�omoǡ| q�M��jXv!�fi�Aɟ��/��z7��&�~p����V5L���-�Fa}	�o���bɋ��18��S'�P�������k�׬��d`��*��I,�u$��<έ�]����e+��J���7�3k��J<��%r��X���p����$�e�⽢Z�6!ɉn9쬶��4]P�b�������7�h\V��q|��·=�D������x��y�ײ���;J@%�С�᭠�,ٸ���ڄN�c����9���țm�/��������N�i&w�i���`���gՖ�y��@��ƛ��á��?8��(�o5V�\5ҩI;%#㳇!��3���GF���}L<�a�q�G!��pE�'������,�D�%�I�z3Zw�hE���X�c#������0���l���#�D�:��BK3L|��!�DR��*|i*����71|��� i�VZ?�'S�Ղ�/V���� t��Y��E�ƚ��#���j$��$�V��2G��~�(g�����-�hU���Ig��������إ�C���_�)6G������o���+�-��p0��xYUx	�x�����XZk�U4@i�ڙvd�6z1�4Q�Y�����#ƐI�~���)9����o!ʭ���.)K�#4��%�_��
�w�H�/�P�,��@n�*���9������,�q������4\ ���S�©����k<x9+IˀґC���3jk���� ����pr�7��g��y�a���ݥ�o�g0�q Gd���u[Kl��*��8�,�q蔑�Q�T��ˍ\"��I;$�H���s���-A����@Ә�!��j�&��5`E���E�D�����_�)%ipp�F�!"0}"E|�3. �V����rp~_3p�C��TE%26e;[��7K����y�ڛw7IocW������C ��~v��J#V���_�W������YBV6~r�k������+����(�&K$#��-R��jNY[�pb)�r(� *�e���C^�zݲB��.�O��-T�::$ ��:������>�3�eYx�6xW��eV�������^�M:��MD��1Mp��e�7�;o/�@S�na74v%D��9����D��x*�P�L�S���l���S�~u3^M�1��Q���Կ)Q���v������sO��-��w��
�t�U[}�5�������:�kX�z#���s�{�&yj$����4b��b��ܴz�%��4�K�B�@�-Eķ���Zr�@KQ���҆��RD����N� U�y�e����z��]������}q�K=�DZ.?/9�VV�z��X&�~9�vۋ����@���0����-��^ �D��P������ɷ@O::Y��~b� �Έ<���oH�\M��HYk�� E�>w�z�"w�·k���LG.�LDL�Z>飦Me����,��|�~�!�5�a��2�- ^�o�ݿ)������������L�t�p-]�m�v��!�Bs*~x���O�PQl��CG�J(Mm�&�\��\�[���`}īt{C��	�;&�0R|�bWO����c0�htwk�PZ�T�\��P�P4��L���ח{q��'��z�њD�{��9hEXI���d��a�ex;��WM�5�`�̖�6�t�_so�j�[����H`T����ͺX�F����k)w�e>����tpѤ΄�(O�����+��]��ȴS�s$v��{�^�q+��uw�x�F�M:2R�"���S���k9x���Ǡ�z�c���%���5E�s�M����}D�n34������`$^U�4��1�(�P_��k�M/��b���!-���w'Xˢ���1�3Y�aĨf�<�p�d���c2Ǝ���"�e�`F�eI�i;��~��h7s$~��ar����e	2��I �55��v�^ <:5�:K�갔-��'AC��--r��D���
 51$� � �{�F˝��ů���s�z���t)Vn]\�����}fk��o��/pm3��VV�i܊��t;3\r��JP�W��u�dϧ���@C�԰�5r9�QNi��Z}r�k�r2��9����[���i�ZH���Ϻ�9~�n�c���c3	azϓ��B�-3og�������+�j�����>�}��g3�(�n�KoC=���ݴ�kn�a�z���V��%�w���5��|;�&����僋�$c��z�!��e�TOc�����7���G.�_Omu~���mm���B����"\�����T����-�WF`5ޤ��Q�=.���D2�~C{c�.�;���:��b�PJ�iE�g�C.�.��;�J�K<�|A��Sf|�To ��!9
r���S�A/��tI<&s�V���&���ӱ��B6]���="�g�J��<�@�iL6�iy`��M��
~m�"<,�V��f��Ygm ������M�����z`&g:
��$�����?�C����rc��ܓl���y��y�V�4�C��x^��m�|��h��1�sR���*!Uo��I5�kj" ����W_zy�	�
���v7�b�>�=�/�Du���+����T���ۿ���Ҭ��)���]����,���i�[)�_dQ�+� Z�T��ifό���ܖ�XE�����T��k,�c�ǿ�������?,k���F��C��_�5 K*���4�ˌ�RG�3.b�H2�S& X������o��
G���`a�*����0@��x˿���!�����������-�2���?�M�7S,Ny���#��춏�R��r<O���ߕ䬚���p���n�g�PR�j?"�d��v�z����HcŽ�QAR�[<�}x[�|��: Q��ܻ��x[9�Y
p%e��(�%�l�8.�G�9�0b���MQ�N�r�o�>{��D�JmLczY1��'�> ��+�7:�>��4�v˰�B���x��N7X:�I(�q���`�K�\0֏�I'�绺bخ�#���?���%n+vǏ4a�.��fS��U���?�mT�iE�$a�8�47�������N����F��;����ᴯL����Y2���߸#`��
�w_p�>>�?+���x1!��������u�l�n�3!�"46#�x*jWFW�~����X�Ku��k�1��qͿ�k��LhQ��nN6ޡ����z����a��k����P�Yo�$�I�ysZ8>8	;��o���e�ܤ�ږs�)�s�W)M�`3n��^!��	�Zi��sc���3�av}�r�k*��+H�wk[,�b[?x�6��p6�*��
E/4�����:D#�A�K������q��[-��P�n�����"P��G�����,��(Dͫ��Ȟ�i_��R�W�i֦�2���E�XD}Ʋ~��D�F6�\h���2�n<f�ޞ�9MSɪ[idj�yE�+1�N����!I��>�x��G�e��*�;���k����gQii�(�j4~�|��Ag_Q�?[.fs���a��ĳ&28�U�f�ኛOK�5?��Io�vv��R�E��o^�h)��/��d�{�k冚>�U�����63@#�1�}>J�4�/?�WS���ͮ]+�/��\���x{t�S�s�$�yB��s��"ݯau�s@��l�W6NN��n��m�⾛_�«r1H*QLp0��ba��;�z�?-�o���ƯO�f���-���?���ډ�5�hoy�9%����V{w�#"O۫�q��A*2($�c�1I�rWv�w�x�������{3V$��k�H_���_�T��?z��=ݘ�I�@2
��;�����>���&�LSSfo��i���Jo1j�#����P��S�Y�w*�����|x�'�h�+�/�+�R��~�[f_�;-��-Ҏ���������ƕ2I]��~~#m�i��v�nk%�د�m�����e����g ���fY��d�Ļپ>2����r��5K�����[.������~�%	#
)zZ�fZ{5�b�T^��V֖b��pH ���oȼ��D�X�oF�T��jxЉ!p2�^��k9ra3E���^�4Y�~2��`��{p���إ%mm�e���?��	�f������#h��f��g�~d5�Ȗ�LϏ�r՗L�����)2�N�)��񜭞�E`aD����m~�c�;�z�?�v��jf�ǝԩP�G��cW}��JƬs���dt��7*�7��`���w�J\���x�)���~N��ӓ�����M箉������˩E���GZ�>FFT �6Z�ݮ��_y�GGz�2I��f���!��� %w�b�Q�P��7pU����d��&Q�&n���`2��O@f��p�e����DC��D�5���OD�g�1�����+��SV�GG��.����8�A,��	�ۋ��[��zӫ#�:NF�RQGGGe8����:n������}�ߜ��?����e�����H���mhÜ@�[�N�_�n%�ޝ?X��NtS��D*�ȸ��o T\����� �o�Ji;�R'VUS3u��l��Wb?
b�OJ3��&~���z�L%���/f'-�0�_F��!_^7n��!�t����R.?�/�$y�fȹ=�~]�.M��U�G�SD!�أ��M;v%?��*��J �Q�QS� ��5\d��H$��]�}�:�%�?�y��-�<@x��s���c�؁��B��3j͏m���\���Z	ږʟ���l⵬k��H|�L�%�c��x�5A��}h�������ʉ:]�J��s
z�p�D~<ͺ��e��M[��:��BEaC_��Q@���P)�&���w��y���%��1��DKS��,E(��h�&���_X�{:�-y�!A����tkcD��b*��"plL~��c��Z�7�.+0���.���Bb<�Wyu��7�A�qAI?���_?���|�c$H�h�x�]��~���l�xX�Q�����B��~��Y�,� V��6�#͏^Sc��%���/�ZC���J˅��j���=��TE�(ޑ"-��z*H��,b�����y���Mz�����e�b6.H�ңdcL�^HKj²F�L�5��ƃ�]/��[M���o�O⪿7�K��9���f�X|������t)Ywi�^"}S��,��"d�uq���t��a!�Ґ�b�\i��&�M�?i��B�ܼ�m	z�Y��ۼe����!�:4�ϴ���^�d+wji�Hf����.���x:�.�tE|���-9����l^������{�v����� �����?5H~~z�^�+���?��k/��`��y��vC<�s������C�6KWVQi�1������G���J�&��h�L:ބK����-�-��I�zL�w2=��D7�/��� mtnW3��P�P3�	���7hhhvw����:ff� Uv�LP��"�25bb�q*jQˀ��V�jОF�k=���4w��~a�~���;$��+�W�aN�\�)��Ĝ|~�&�m��7Vz=���I���K;v�W�o��
7qi��Ŀ�{�͙qE��>/D���af�j�l��Z.��_����T^Pm��37`�P{C��}�������FI%T�L�m�����l�䵶v���Ա��Bc�hĎ�~`����*��@L����6�QQ��!��3H��\���5��S�P�԰l�spx��v�� ��Ll�X"���p�Im�&��������8e�	7t����v�ł�e�:�"��@������́� ���P�.��!�*�q�`yc/�Γߩ� z��A���K�B��t]��7/O���n��O��2�)�%uL��V���.R:���F"ΐ̿���|'KqS9C_�H��6Oϑz����C�J�㢉���:�o�[=������\N����a���n��k�%ԊB�r��ףݐ���o�f�v`]�$�u��Y��$�F���I� �#��H���XG��<�)5��y�@�v?�mҹ��D
�N����3���B�*�����dϧ�-�-�1ҧ3�z��9~VV��mQTU5.��q�R3Z�ˢ��UK�Q9qqT���Γ�y��V�>�k�-3k�[��1�;��n��f�g=/p��[�^m��TM
��,YO�����0k-�uE{�Q'+���@F1���ɬ]�'s�����Q(�F��`�^},���f,�V�Y�z���&ƳŌRm3�Ums��Q��,;�bn����m+N
X�f8O���8ӌ�ͳ�!Ɗ�/�:�W�ג�w��<��P�jߖ+\ﵟX��U�l%�J��n �������7���G�[��~T�\(�&�N>�u��\��S��^�Iq�£4�_#6Ȉk�W� �=ڌ��ǒ��ya�h��>��B9"��J�PL��<�	 ��2[o���^M���GCn�ċ_5
	�ksRg~U-K��_\�W	�dȶX $�y\�&h����N���Y ��n�v;o�%ux\[G ��I�瓤��N,Z�m�� A��|{_��jC��ZG�^T
���D��e.�`q%��
���h'Tk�_�"?�0�rդ�=Bd��9�m�1|}�'9jU*d����8@.��qW����?�B�kGN���u1���Px�?ؔ��0YI�{)koan^`���o�e�3ۡwW��-�~��߀� ��AG&����V`��I�.8If@��I��<���s(�◣��X��]��a�����7���P�w?~�XK�j��t�����Ω�n��93W��6ǾQ�.�۵W	���.��-V�K�-9�00����"��s��x�C���]2>�[��ͼ��)I����Q#��-A�^]������
��J�Y��ۼ�Y1�٠x_��X�,BrUDU���!�p���k���i%�H$,��=��,n'	1+�������PQCp��I]]���W3@� a��>���0n�D��ʉ,1���-��qCj�wu�^X��5�^����,��~C.��7��ú�o�A`9�g����1�}�F�%���ˏ�tZv{�$�TUy��g��?Е��7�	��E���gy�v��'�տ7��_q�AI�G11��>�͙c5�4�5������)�u��l,�"�D������b�{	�]v����Y�;�y&��{d����^�	��{��j6��*��.'9kxɊ��
8Zơ��h�`S{�m{�;
�E;��Xx�4�F���>G�Ӣh��{?p������n�^�G׾�W̯�/���p�ll��Y��'�:� ���gT���,��e+iW����f�w43��|b8�^'��N|��9!X(����Ծ[��Ӎ��܏T�yC��Z}�`���R�Gw��x�q&'YD*9�d�̥����opc�{�����ٝA��ʭs�.z��Y�r�<U�\�럇�xxF��g��n���k���o'�L�b���`��y�Z#�P���E;R��Z����aP�c�W�B��Ph}�m��>�ڝ{�!��Ɔ����6������	�޽�򪫕onli|w�⏫~g�1�3,�#FW�L�{r��tnuAr�lXʏ�M���u#���3F��~f����f��`���7��K���;�ߚ]���C����O+�z������� �8u�xc���Uc��R	�l���hW]���l��;��j_�I;<��a���I�`ʠ-�y����pں�%�q��ļ}��{�g�:;����9熪�Կ|1�A�&8_k�@�Bh\��P�V�:��{Mۯt2�iU��v�w���,��(��\Ri+��~v	�SG4�J��-`R��	�����]ն旝r��;Ocj�2W�ObG�z�Z�lh��.ɯ�P@2���׿学ԧ$M�����ۺ#s����C�F��I���NZ��6(h���6x���s�i]X��~�2Z�`U�+�,0y��5��m�l�|<�6���"N)U��H�?4����șc��u�������R�l���]�ź��ރ��б|���7��:vk��m��0�T�Q��y���&C���� (:���-K�j%�PW(�v���ۣ�jܝ�o�;�.�>	��L(�4z�x�[#�J&4�G�����ɜ��}���Pu���\��M�.�����e\K��
�Kxy��8�Ɉ]�!��q��RB�#��x�]�������s]A��'m@��`�� ����p���̿�ڭ}������(�(gk^PSg��7]~������5^e��h�(�.���JY�ݹY�zo��	q���y�s��-D� 2�R4�!K܄jz�|B�W����W>222vP"��r1ֽ�}u8��Y��Aj�������% 7�51���*毴�׶�U*�+�-_#B�eׯ#l4V4�4�_Q�s?ּ����j��g��s-����Y��=�p n�3� ��Y�I�Vz�%�Z�������^���|#A<ߩ)l�>�s��g)j�P�ܰ�����&��4?��?�r�/#S��>[�����
���5I�Z���t��������;�<r��w��#@yꎳ��w�I�K�}�T��k��>w�m7��'}�:� ���hXhYk1�כ-st�V�ش�K�XJ��ҭH��S�u��E�ZL-ϐ�=�5E�q�$�#��Kc�["|�Y�p��F+u���)���)�q]��w�x�̧J,��,>s[q�*�z�m����yI�j���r���s4詄��p�� 6*iߋ��V\R.�����0aj�	䥠�#S�Ma�(Ĥ�'���0u�h�i�i����u`1�5�ԍ9�s�.���v�C�t��v���g��t}Dd]?�T�w��]��{��@u����ZJ��}ȶ�<�Y/S��0���@[�!2�˧�7�<=��"���1�P,�%f�rHL�.���'囗�>���q��u�O$RPV��c�T����t/eQ��"�Ъ�Ҕ��ɂ�_	ǩz��1+w��,(R��L�G��,�Q��7�2���)�Mv��� ��!�'����w��O�Џ#�b�(t�r_<~��s���3Z�j���z�M�8�ֲ����.?
>�nSԫ�ok�ds	I�{���s�8���WM}���q�L�r��*�G�ƀ�"N�w����WN�M�F�JP5V��V�̃s�v�^^$�aʒ�˓�p��@�0�QL/�,�������ː�h"�[Zm��hN�ۭ7
w�{���i���թ��	�O�!�_2Վ�y����B^Z����[LٯI���W�(�]?J�ɕ�^g�v�EG�v��i>sC��[�R�Wr0Vs�ʞQD�*a�0�ı.f�a�UB����\�A(B�m�вݠ��b��|h��q��s	]QJ��HΩ�e�t���t!<�����f���`CO!��,9���oH��>�-;�[��
�eEٚ��3��5�ب��Tux��k����?`"�ݨe�.����Mb1�L#j"B��7�+?�����q2���My�w� 0����/<�4;u��>;�d�a߬x���Q>���걞fY���������J�)#ݣ�A�x�'��0�a�t�V���G����'n�����w�x�q
�ە��d#O������ߝ�m��<�"�8/�_�@��u�x��],D�����coF�=�����Le�"+^�?oD���m}C�z�W�1�K���!�@Ϻ+6l+����P(���I`?���K�ͬ��u���,q����1o��]��' ����@��3��%�U~!��B����\{`0
BW8��[o8���QmQww����a|�;PfZ�W��8�@A1������h $<���DC��<+2}���kh�N�<5����4
��d�P���H�T�]�Zq����C k�J�� ����f9��z���w�JU�t��-�~ �ӕ		�z�5(&�K�[����BP޴C�#9�L2�z�xx��BQ�{�Hg�X��� ޢ��8O��7V�d/����:���Q`g�`^�����=��A#�T��0���mՃ�!]�'b'}���U]�fީIO�s���Q�KRc����s2�U�Aʯ��}�'"��<���"#���z_o��WEb��C3�pť��M���J,)��P��XK;��Sl3f�6�J�PH+p�<�cp����{�Y�7$�u4@=ojյ��h�҂�N9!�k����ݡqzӕ�T�]�-��3��튲�T�3-j�����a�,�K�������t������KG6���X�� k���p�b6ƀ�sR�ˬ���z�V]��K��6#��ф���x�M�Y�����
�3m������Y��=�TH]���y�څ�d�2=�4�ғ��6�fD�~hWⓉ+�%�(k'�4^m�%M��D6�\a���0��	d�N�J��k͑$g�X5
�ݞ=���-�T>t��ǩ�����4��_-@�ɇ��
�Ƌ<��6� �n����G��G�B�PP���W�ܞw[�S<����q<+<5FX�H�����E|w���9��ef��!>������-Zޗǋ��n���GZ�5_�� �Ʀy��:�!�����C>�X^	�;Zx�%u	pB@��D�yi6�X.ő� 1�s�Pr~������0�?�v��-�p�c?��=����^4"#�`�0�<ã+�:����k��_���])�qb�5�O�䕆��0����hj�{iT
�{�n�1�o�;��G~�`���C���p�~����P-v|��jQ�҃�DM���@�=�1F�~�q����fw�Zw�i�[z��5)]�7��y��3N��)��E���#ꭣ����q@:�� "�ҍ�tJ��tץ�A�����N�KHww�����~�\ֺ뜽��<�̳g>��!zz8.RZFw
ؚ���=l�S�=~�ؤ���ViU�o�(��[����Z�g���65���ھ�?c����֨i�$;���K�����WDxڷ�]`�<W!i��[��o�o��9S�q;�P�0)�Wz�#��j�#���YA��$a��0b���M�{E"6���&K��Y��t/��1W�tɗ�FbU%�����)�C�,u`���
=>������o�)F��cKz�ڰ�ȶ��d�	�g \��� _�]�n��X:��J�����_�)+tc����S�ɪ����Ah�x���dg���]`��R�1�� �B�G�F�������T��0�w/U��g�|p���,
��b������`� 益��\��7S5TK��QȂ$�>����D�Z�ϻ�Q�a	>�ɳ���E�i�}��'����%fWa��,{����`w�(kDv���	�K7�Ph���޽���A�^�%��,3���6UA��Q����^p��ڞ����L�iJ�j���Ep�@~�A�%q�~�Ulls�7��u��t�T�(^���@x�Ӏ�3�:�nz��`�o�@���٩�����P�(�NM��3�\���L UpvfE�A�i�5����sVK�@��e����0��;�I���g���=We9�U ���8S�Y	��X�/5�'�V_q�p�v�L�|Z5:��s�¾;0��8x��~K�����y���Y�����]���V������?u�\����@���������6Q��w>R��\�x��\O��J�iڻz��k[���0����E��?E����W7�T�2K�F��cN"Y�C�%�\2�Y/�^����Q��UH��1s��i�?�~-z��E�{���w��*`�l�W�_����.7Kl��B��J=Ijj����|���Ǝ�ǖ�������ɘJ��@�U���N�p���d�ˉu
z-F)d�v�{��c���F?U"5�c�wZ��1~^nL��#B����(�V�T��:bOp�fdg�-�[� �0>Y��ip�l�������
���$���}P~M���*��d>��C� ��K9Vi$��\kS��6c��q�A{���&��ǜ��<�e6�މ�ы.�ĥwgV�t銲��GaFҭ��=$�i-	�+�+1��p��R�>ެ�oɟ:�8מ���F����l~t��?�}7I�����kv��p����x�4��a�|�c���{FOI��h�����%,��S�gKGr|�x�m�me���W����h��?=+��j�t�&�{f�}��B���0Qz���'*�EuI8i�f
C����0���%���j���L�>lĈ+��@�xS�'�
&|;���5Cy�9�+:>.�2z���w�=Na	�K��;PDv�9��_�E��z'������E�O!����.y)�`��B�~� R����E��ܠ���D�\�3�e��}a
l}�$��C��f �]�R����=�����ԯF0cv3R	�_&7u�]���Ven��Wp�찒�<�W��:stKR՜���C}Z��$��Wz����v?��E���_��?u�}�|9Ϛ�!��O�׶��Mnz=E�;u6���ֱ�;컨ٳB )3�S1���|�Z��ˣc8K�2i�e�k�o�&�'����ir��oS�}�lF���`�ɀ�a�2w�`�}�VR������jة�w�W�m.��a�>�o�R �;;>!�d��+Y�_$""�����F��_�P�x���P�L�-���kQQQ�k����c6²b���jf� �V�/��ퟛ}8z�j;OF��b�7�cX����������%�1���;���ВXO�A�1�mZ�������׼�1b�6�}�M�|��9��6�I��0`�>��W�BYNm�p���HE��l����i댒�Q�O��*"i�Ob��|��k�����������Pii��ь�
l��e|f��	�J�Ji
7"���|��(~(����UC����܈��������E�����e`��
��^Pцr��	�{�q| mp���m)����a>�U�t�~ӱ)�
|7VPLd���K�E�������CV�(.$w���>�U�@s��H)e���$�a*;$���N�	�%��^
�rh)Ƒ�g(�����@�����z��i?��ؘqѡ���1����֙3F_+�n�lti���]�=DCMm��I< v0}�R)�\{|���?5�4�C�qؒ.���'S<��ܘJ�N�]���cE���2F�]�s<���^W��H
FTL�\k�	���,�|��+��$� K���mi1B�ii~>�Pr�뺂�$pf��G6���A�iȬ�FJ
�T+��`�n��vzMU&")���/�\���L��#�Jd���o���<�ҷ;�!y�<D"ya�'��T�qC�&����C�bF3�����&+����S�G���~�!�/�h�H�,�$����Z��|�kz_����iX;��b��&�ƪ'E�=��x�4��eV	U.��mQ��̗�u3��K����=9m��ߔ1�Z�p
�4(��f�Y[s��`�X�h��-/\�Ea�jq�� ���4�]`�S�k�M�?f�Y#Ѵ���i<g=��%1z��|,>Vk��X�P�>�@��hAj� ���b�G�U�������ƒ�9��ׯW��.��γ�w�������Ҫ��hR���P�\BBB�����o��&&Vu����`X H���z[�]���^���}5j^��8����|��U����M�ý���8&���5�Cw�Y�8#F?7I�7.�1DXIQښn��Gy�4�]���~ge�S둌����(��"����U?��b�����9�4��&j!��nu�[V}4	�$J���_H�H́���es��8�l��<�17	TI���[[[�}PN�䢟A,�MU �K��$>��D�׳���)@��~��d��R��VY��*S��͠��2ER��Ҽ����9��\�D�u��n�̎�?A5�k+%+�/G_���K���a�/�L�c���⠳R���GU�;�ýB9I� HUW�����<'� @F�����*�������Px¥�ځ:�՗wW�<3�A'k�o3���c�̜���ol.pjFC�oC?GT�.��L��z���^�=86\�a�W�{uE&"n�X#�8��9�H߄q�5�=F��ڳ�~���]�a]�E���z����)$	��X���7P�����g6Rw(�x�\,�av���xR]�� �o��
D� ����+@�*�H�3�_��kp�˜x]�G��RӬQ��s�p�hr�{UC����AU��~��d�wKk�����m�K2��s;�o�>��|�#��6|�nUg�iv���@�'C�<���Gg���d��j�n���]M*��iϼ�apĮ��f��}�t�
Q�ZA%��b#������}��0��׹�kc��>�V]x����*�������ժ�m�ݖ^S[�K����丫� ڲ!k+8=|��*�Ę�:�9��3����H1e��$C��8�8�q��f����?��*F��پ/������ջ~��]C�����c��S}���2\Ҡ"�bSF3�5���DE���>�-��	;n4�ݭa�eV��^�n��5�V%D�9��� r�|�M��Zfw�Y�N��']�:)�+���y�Ar1���;I���E���9+ƛ��(�z�
����!a��e����n���=u���cg���jwd�ò�_�n7YЃms�{PG��G�qs��Gr�ˎW�<�ʏ�����£*�_r��Լ�ڻ���2 ��Q��Cp���!�&$H�g*���
9jW!���Լ�b��+Y�
zuU.F Lk:�<4���&����e�6��g�	�}^O�j��`*)Cc��.YQo�����2����}�OoKqh)�����۸n(�;�ջ@�~v�\gE6����Z�\��us� �����q|D[���?��Y��o��r��<ρ:��fqG����e,� �	LH�q�g��-B$����k�o�<J4:ƨ̡�nʴ5�b�!�m��ݝ,�}���e+ßBY�1�\T>)	�n�5bj�;!r�/-���t��:�^�|�����e
,g)k�{2ތ !q%�L`ECA�	y�#-�Ul��®M��̈E�V�x��
�{��u���\��jW�4ݤ4��l,>a	b�DP�j�?��v`��i�����a�^L%�;	b���Q�ӚX:��Z� �D��/�Ò�Ҷ��99��U�L���D�eK��g��܆�!��!Pk1�mX<���p7�k%jj\\0Ĳ��
�������������Y��*)Q�;�\�� ��旰�*�9�q� v}̢o��y�6l�Xv����jF������]g,��U~��V��bcq��9�iz��]�]�Tn��N�wȼ�
M�R�i�9V�s�dΦ�\/ߗ�u6��허���+��Vt� �,��%��вM�]⎻���G�[�ʹe�Iܖ`r�+�A�
?��'��[��y�<�]�B�[�ފmD�IX�-o�-����~�4���2fFO�3NOWf�5�lU/�N-*����?/�Ő��A,$H�Qp7��10���I�c�}�GQ=�Pʬ����][W�z��!��PM.������ʙXx������9ˌ���Ē�V�!妖h�nY;}��>:�â�;����d����fd���QӤgͳO��Y&GlY�-'�C��$���7�8\6�N��<WB���݀)���&&�`�l�.�D��Qf�Ƣ��OWB�d�o0*��3k�K��A:��`8Q��n��^ ǭ�� x���O%a+uZ[�*�z1.#�]{/"@�G�hĀog��n���G�OJ�������R�>F����A:_C���<o�"y��5D��5N��7M�0����c �po+��8d�����,e��X��A�yϩn�@"U��F�� ������:_���z�������<�De')����f�=�>֬�e��W�#��#i��.��Q�ߤ�Q�tϚ�l�O���T*̏L��\S�ԉ�~\�Fh;-	Iօ�c�qp��G<Ǩ����"�g��52�蝖nF��w.>�li��U�
��������9��wn�	zm\?��H������ߜ�`����O�m���|^3-��L��Fh����{��'�(6D�r��� T���s��4'��<{v��q��)�6_�e��<<_�pE�Z��7xm�z�[�m/Zq��\i�/�Z���:��ۚ���g߽�$f����F�4�1��Wթ�'��w�?��0���r�/�ǡ�b
/���ql����=�%X�ݐ����j ��|Ps�Je�#��;�Ɛ9�`2���R[�)�tm;Qo����~]�4�K�K��eA�E��F�-_���3�{ktؓ�����/W<���	g������an�De� a�n�fJ�v:����3�,�	�
��;�e�����~\p��K�a1�cyL1$& 7E��ވ��b�@/"��&Wg�D*�����t�k�}{E|]��*ŷ,r�l�\W�H��Yq��s����q#N<<<�s�~�7g[`9��tcp���B�b���氤�9ܖ/��	�TH���a+W��*��I,�a�Y���텣�KY�֣~��"���&�9��(h��#W�R�+�.��Q^c�b�H1�8��tAf2!%L���9���R���"�Y�;��+2�r�4Y<0�Wʜ�߷xP	�h����T8�����D��U���>�^��<�
>�� FTe9���*\����7	��%~���`�A��jwߨ皵gQ�tP����m��fq�,�Z��xA5X��UX���[���+�����c��>�90R�,��,�D<��u9&���ѣ!ٜ�H{Y���A�����>yzt����p��^� �c�J��� W���+�?���Y�1}���s��Ou*�����CG�y��y(\����[q����
���⦛�,��)�Ex�����I�F����x�q+Nu*L�jX	��4.��ٱ�Q��U`k_~��{��u �J�,,]��p ������ϯ|q����>�y)�k�����m�s�"ˤ}M�"�,&�;�
��,%($��y��g��,�?[NMz��3OM�8kE*�a�NI�Q'I��8�P���אE��
�&�tm��(L�
&Bg쯹�V���		6z�#��T���ޯ�")�_p����	%Ѩ��u��N�����|8��h�ݛ+��*aN�j�/wB���5Н"�r��ؤA*�O$��)�`����(` ���
*@6���}ç��y3ב�}��%is2���Y���s�����5m��9��F ���᲻�u�xj���o�EHct0���!�
�U�ڌ�
e�NL�P�r���D��=J,Q1ҳ�2P3���XA� �/�03��֗�E��!$e�9��[?w�p�0w�
 �z(Id3�� �uX_������w���3�M�nG*�d
{�Lu%ŷ�%ă�|��!��:-&�R6�/������5����LÍDF$�߬�d��k��N8���\a2��HW�m��H1��㕮_Q��j|{)��KPC�f��k6�Z'k�`�7Z�Æ-��P,�݂���#�t��$!��G˔ �_�[qo<���I�_�΀�h����;fl��Qi�&F`�PW_�ih֘�+��]����Aٽ��2ϒ#�$�F�P4�w�g\�R7�z�K[�)�8����Fv�"6Y�o&W�s-Q�l$�
��-����>o�GT��ſ���趤��L����u�N�%�S�u�~��]���N��L �V?[��:��R��s�$R����'�2�y���)�d2Э��#�'����`�N����E�*x� J����6�aར�U�s$���|8a��G
o�G3��nFS+4P�"�(Y.���Ė�C|�u��vGW*�rGS�C�ً���F�v5NY�=����t�=��
,f�R��� ���Nxv27`+�y��"��o�P�
���HǤz&�f!]'S��>ajv�$�4/��#�	,�y��[���hVP�7
>�iV�q<]�R'0e��K�$��f���w��_��FV��x��r�(Lj%����!E�/?=,�9PhY�S����;0P��������1s�=�Lv�T2�o^��h�I>p��ٲ���7��-��
Lm�h��S,�9��=��s�Iɖv�� ���jͪ��M�:s���*�B6�'y��W��o�K���p�
���$�`\i�ؗ�����A���t�>���$�v�m���������*�y?�A0��	�do	�J�>�|[���� ����}!�{���&��'�z;�$*��~֋-��hn���&��y�����>8ѻMC@� n����� ��ӁLL冞7�y���@J��3�T�ߔy��O�S��
Y���Ʈ05�J�ɀ�n�:e��qH�����:w�zp��G��w~�҄����|Gf��] {�<�U�7�45	,Fӣ��#N���2���������"g�R�ru��n��E6��m 5Q��%;h�9n,6H��fƩ�j�ۑ��v�Uճ�#�v�+�Hݓ`$�	�Ǚ7P।���vw\�Xr�-�)�=59���Ȼ9�Id�	����Z�˺�����^ as �nMIkkSrVx�x��(�y}QFo�j<ﶽA&���Ju�$S�����7����۰��A��2�/��pw_S�@=Mk^���5���2eT�}��@����:,��,�zc}��	�f�f�T/ܿ^a���r4I��|s��T��?]8~��el��S���p\hp���;�r��߰*�r6F��,e��7-�v�ڤ~�ԃ�����2�WݴZ���\_�l�/�p��-m�a��)�5�7��ؼ����F��w��j�d�U=�*��Ab���;��Z�	b�ύxÜ�~<B"�sRs_
�T�����}пhjj��3�?W^ic1��wu�^��&��S�����O���ah��ە�:��U;h�x����nFnU�e������߾�$�|��4	#���!��M.�����i���Z%�
��>O\�D޸#K�&3��t�%P���k�=M�Q�����Zѱ_܄�Bg�CC}��|��|�T ���,�F�������X��)Yn��f���`j��a���v�_غ�� lJ�� �WG_�,���� ���Y��3�TDn�t	6|ߙ�l�mْeҶ��x��G���WU/���<Q���������2@F�(��y���r�ߢ�Ҏ˳�o(4�g��!����¢%]�Ȱ�1^��1��⧟�p��)m@]�����ѵNlQ�����\=X� �8ؒ ���<R=T;��"�ˬĘHXM����5R�3��¡��@Y�i�NM޳�SZ����D��j��S��I���(��1<��C��[��v�+��"tL���
�u���F�(�m̻_z�Qc�a�^m�L.ΰԶN�~u/��,^bĂ*�4Ψ��oI�RG,�����{���Hr�dhr��u'$��p)+4�P�%��jz��9�&�S�!���XA�Ʃ��D�|��}E(#�{*e�}B�^�e)wE��ƺ9DS����)-:�/��6Q(+&��i�'"ۍ	/��
�F6
Q ̟M�a���C'T�F,�q�Igp����~�S�[��M�@x��{~�Ł�mrs��J@�g#h�CW8�O{��j��&��r��*�����ޢCó�/߀Y�{ȼd�J�qc�Oc���w�4��u*J�����n�a��!�A~�z�Qt}"Yf��;Q�PD���j��c�	��p�:z�vW��)��J�|a�=r����,���tm�E��?X�ykO��*u0ʡ�F^�<2�}bAw`�#�E�Y;5����сQ���R��g�9�}{�U4`��$��������Kv�|�:�s�$s�Χ�ۤ��Y�֣��:�ڰ+�_��gX�Q� ��T�J���I}D��᯶�9���H\�ѵƄ[�N�^+@�V3�&���ƙ���*ճܫT�f8� V�i���Ov�Z�z�t9�B�`����.LW�>'�
Ŧ|N�M��W�Ķ��>�4~ɝ�=@>��Fi'*$���c���:�w�p�%�7&j��8�(Oh���/�:18�!z�:��a<��0>�;�a�#!�WU��P�?2������r�i]���n��`��K���"������>�<5q���#x��L��f�y��A(�=���"�������P0�	��\\\�}�ƚ�p7��$�)2�r�[Ը���~a;M���B�� 9����S-��Wu�ce�s;�O��o0���kM���/l��Z��G�_Ù�K0����X̥�i��[H0��Cg�H�AN�q۷U�n\)0@ ΄�7řs��k��өw�6�9�c ���lpն�`�_�W�b�G��	��;����
�*ݑ�����Y��?'�a��Q��-��J����	?vLC+�-�_mb;a����JD|������S�a����c����ή��M{���������oiM~�H�%���"Q�Q�Y�(s��.�G�G>�)��ڶ9"�4;�>FCX�i]���2[��A�5�@�~����v�2z�2��Zc \�	+)�E�����C��of��A�b��f��)c%@��S�1+הoy̶�RrYe�������V��5����{PO&���Ʃ�E�C x�W�G-T핧��f��c�� 6z�qb��9IG��yR[�Gx&�@���<ׯ쬬�.��/)�����3�2C���������, �����	)�������\�Ww��>��Ԋ$�u��Fc���P��������u�V.�e7.��.�-����u-c�42��H��k���X�:�;� @g$R\����L�����ӭ��C����W�a��N�j^�^!Qv�V8�G���L��e�����m�x9��9��Ф�0뇆�d�P�ƈ�F��8��!V)__apѯ��)����mo�W"߸#4�(�>���]�f�����ݚZ����Y>E�
/��xӇo�� ��y���2��\�^����_�8��	���C���qK�%j�*0��P�U^f�`��n��5z��4�_}�snఞd�����乆ŢW�)�q�c���AN���33`C�X��/=.]t���.����y�����f?��LB��x�c#ݧ�z�#��������R?;�N4���Y��'��EO���%�+\wt~8���JD��~ʢRw�4F#9U��C�Vֿ=�����s����5،߆Vz0P���R1T�n1!v�6Xʈ����}فkL[�bCE �ρZ��Fvph��`����1���9(`UJ��"��W
8b�:o}���%����W6��?�H�`f�b)	&t�ϟ����P�j�&,�Y	|���+q��S*zp�kʟ��6G�Z	fA��y���+�4F	f��ψϚ+�j��|���Ls��IV,Sk��e�͎S�ڠ��s+ͣ�v��ب������Z���2�h�-- 惫dV���#�fdv�b��X��y��i�VW�J�ѯ^��c�N�p�c�2���ee4�լz(^�va�D��ED�i��Ӵt�/B�:]{V���y�eo��z8T�-�L��=G��B�@>��s3�>�љ���-�[�7�(^zv��G�x��h��,:�pg�Ý��/7�Fo�;l<�@��B��E��tw� ��Q`�7�~��l�4�4 8y:�i����2C[��V.Wٚˋǣ���o�!�� C���=6�u��#��ы������֒�)�J�]��ޘf\��"F�Q.�v�.w�2w�:�9�:[yMg5O��k�- ������L�.��B'�Ee�h �2ddc�	F�g��������z1�Ü�]��5N:����`c$��"	Wp2�k�}&�I�.&칺���6U���T�w�"�w�`y�AI:�t�[y��� H��ҽ��m�=���e�Ne�v̿����j��)�,�B6�(��&i�5���$�k̦g}�)�>�Z�%��������.��!�'�Z۹�$#?��s��do��'0p�%���;��c">EfJHs��̏�>LYJ�~�d�h�ńjIA�s���� ʬ��\�*l��3�_�K�mc�<ۤ��D��o?g�cr)m�[�!XM��\2�	d�DH�jR?'�
'i4�=`q�Ͷ�
�s�}�4��`D|��x�����}���'z�H�(���C /HĽz�q��g�¬w�~ܧh�N�k ���]��
O1�`�Ʀ����IզQ�L�c�=��X��'�{��v8�O@8��S�5�\j��Lį����!_�������'+�C[�Ow��a�'yu���Rqu���u�4D�Y� � �c
� ������1c�L��6��u���sjk	떼�K�/߃�j�Zn����|eq^�;i08bƀm��#TUT�\�����*�O�\�'I�	ͺ����c��1��r!0,���!�N���� � mD�����|�����M�g������E�������`S��v�Ě�x����E�8X�)8��łEٹU.����� c(w�RۇXYY�M�譕* �JIS����XB��k4�T'd8h��`���o~�?̸��CJ��W�_Z(E�E	���Xc���e޺yI���r�B*�?G�J���^�t�*יY�R��Z�F�V=���r�d/j-p�]��{\S���1�1�+�xNo�Mw*�"#��.H��C\\��>4T%MR��YF���R�s�Yp�:��VU�Ȓp[dVT�i�t0�56C��m�
������������y�ݻ�Vm��FmI�.ڷr~<3��d��ъ�X���B^|w/����#~��]6�U���>��qܗ��KZx2��@����c�jw���޵���{�YX̝��%b��x�i�p1?�-��^��3�Q_*��)������CJ��\.���`�w�@
������Z/�An"z���qhA�|�7Yk<�Y���q�k�|�S�ԔyUl�J��l ��M�ܲ~�ᯡ�~ĕ�����_ ��
��p @������x�Wǉ`�L ��y����(cɣ�&�+kmބݰE�8D�@ԀLƾ�o<H���pꇅ�b����$�M4����|�ڛ��3F_�I�YY�{�%�66��Η���s���opr�~�]���1�<���#�� ;"Xx������H�R�:�����F$��c�/���..z_�D���`펃(7\���VWCEL*3B88$��!~�_&� ��_�c�� ���!܄�KRYY]�g?X�����)u�p�/sZ���a�������9_E$��PL$di�K�`��é�R��U�\Cq� ���^��śƯ�5��{�F$|u�5Ҍ�NL����ӝ�:愎�%�I�DYݔ_��p�<�lŌY�������\�u;�`
ͥ��(۷��&�|�)��]f�{c9�{oBB�Z���f�:��_�٤~}�����d�F��;[a�t��
���P���r� ��	�-�9�?����=c�W:��(L͗n���մ�3�\���tG���ś`3�E,~VL �'�;gg���d<żԵv�JT4���+��u����R�>���!��#_���;;��&0���5a�����\p$���̀����<`�9�^�D��s��z�:A=��,�e�������%64�V�)S��|/�Q��x�b��`���9��5�Yi'\m�-:���U������1��］n�	l�	Zb��&�du��������dfE5��+x�Ӆ[�H�g��������(��La�u�:��=�噧����4ع�׻�����C(
6�O#Y�����bu����HD1���>=�Y���`-�������!~S����:�S�%�@��&��2E"6��Y1���5�5�ru����v$z�u7�[�rMCAa�-��2��R[Gmt튞+�z��4q��	�E$q�HM�L�O���Z���#�����T�T�~��]��;����`"x$��z��1�nُp@��ݘ��%��444���9����F��� �ɮ!����n��8���0�Uɰ�]��������h��}������U!����K6��~k�9����S�2B��e��P��£�����:U<��N������Jy�����|��-"��F*�|��"YΊ�t!���t�������*M>X�\�i�g��"�����/ɴFs����0�9��n�'+a���L	��v�t������j���񜷝���s����{6v6��oz��L0wW�^u[����S>��c��h��Y�s�����~P��Yu����9%���6�Y�l�<�g�膳.F)��i-j�Z1��eyL� ���@M*Y� �~:S丠�Q%����]
�J�R�Cӧ�0�N�l����ޡW�����E�CBB��'��g#BG�Tu_���W)��ފ���%i��
/V�^�ޅiW8οw�&'}h�"ߖ��Н�2��?n��GC�y��Jl��*�`W���v��#��ga� �C=��ټ�/H]��P����|�����^���B�W�g/�D�G}Ԩ�H^͊��L`Xg˹@��T����z)� r00��a��J|��%i�2�lx�j��E`�^{l1��}����ډ1�ܜ����YS>]�������d�z�Cp̥ d�RD;	6�a`eE��>��xF4��]=�$Ur �z���v���#��H �Y	j����^�?%��)����;����?L�K�Z�5��Ϯ��d��	����G��� i���$����WR�	:�3cp%b!}K簅��!2�g�Æ�/y�_�P��8R!?'O���F�k�����}�h�&n�������*Ҡ"���`��PJ�|y�E������ŝ="BB�'�]|%�# ���3����o���-��D�\���a��/�)�[)�كM0>hu�O_*V�ǻ�Jt�����_m!�f�Q�u���:J��NR�����\�1K��	Y���Zz�A��:��9޿`�Ͷ;� V�U5�Q�U���¤!��ώL&)�]�6��=}�X'��=m��qpWtr��4Nk=+�0�N�C+�iŬ3��AX�3��ҹ��og*DQ�h�;�=�������C C�A-�`4��*>'ܿ�p#�;�$	�M����+b��lJP#�N�������sC[�\�xv5�([K^f��%����9�Yx�F��븂_���܇Wh^T,������ld��`�3^�,%,��sٰa�����UI��pX������S���t,����H��B�H˽/���P���) ��N!���LW��0���O����i��Ɯ�>L,w�-�ʈ�p?�<EQr$nG���{ɘ�;��^mŮQ
(�X/�����+' ���M��Q�������لs�>��憎���tn��:k]�4��/���>�YEƮWI�^C�\�R��Jv$[�4�A��ݥ	�=�J��R��S���ڷ�t9$^9����c����B��G[CF3� v�T��l(.ao}4��P�G)�����J�8�u�]�����F��,�aL�<��>�{@yy-0�:%�@�P<�B������agAb�V��$*����C&�9q�YrY2W�Ϛ?^y�s����x�(@�ܑ�]���?r2��B̥3�`WOs�goD5���bs��<&�>��R�pP�2Pe�G����pG�純���.=�_kZ�^�D�@/S�Ⱦ���g�{��o��s��B���ÒBh�������֒Ȗ���@̂_:}�: -�$�A)�o�VE/E'`��Di(T��2��ϯw`KhUmm*O�������ꛜU�D�g�ӈ�t3�(<�P��r���+�D �y��b�Z �7�z2�K�+l4�@���i�+���%�+Z'��EG�f���P��o�h =��&��Y�'�ޓ��$�q��fv���2��,�	�39�ً˨�
���ٚ=�,:{a���������:�����
x9 =u�+����D�"�X"e������[ߩ���t�����n�+�p:x�wA�dy��ј��e[S�M"���8>s�Iz�&���ύq�ɳ�2�3�!�g����[+	�yN�+���xů�#�������ƻ[�(�{�^�.$��/^�_�xE��pN�f�U����+��{�z�)�M���u���S��V<�*|I
;������H���'hmO�=�r�����$�޷�ς��qO�t��J{Ӎg?x�����9����s1��0�LT}��R���~7ˍ�~��������	N��8x�2=N����<�<�p>k�)�S(-!q9#�<�׺��m�hB�c���g��*Kt�,�?��ͳ�E�Me�뤧H�M�3,�hͭ�=ؘ�,(�}�[ׄ�ܪdD���oKן��r
D��5��
5=H��Q�ӋN�[�d��N��@�����d�y�ls1v�����|��b��ڢ>�
s7�q�|�;�3Ɠ��'��i-5�$>��j����=���$t�_���l���Nͥ���b��}�1f��4/�*	��ċ��\=7_*�GXf8�bd�~9��Do����^��a�yL�����d�'�MH6�j��H;8g U&���BZ������L�O�D�zZE��{������q�G��$R�2u���Z\��Ŧ* �"!$)9ހ--8�|�z��({��b9����Ho���̍G�箳�
��)��~��fs��_[��@�t%ɷv�рQ)����	��h$WJ<+=K�C_�x�0[�j�%��<\�<�z�?�-Rͺ��]R��
�?���]��*�2�繽���m��*�)2z����+8���`=N���3�!�*�A�1l��\��8)|2ff�pвяK%u[���E�R��g���%nˡN�e6��勌��X���ݕ�8%JP�!s�|k��}���78��Y�=f�4>CI�	J��&�7э�J��P��<������4�D�Nn^5�Ҁ$�fK����"A�{�lM�/H��Ӟ�.����;;�`�*�QSX�8|��W���1�%0Yzrj�`�����"�B"�fS蟃�5�J��!r���53"}�4FV.M˅�%�`�fJ	�L1zP'�V�Sa��wVdUy.���7�0�'�Qؔo�\�bM�i'_��we���8��;two�T{�����5:�z\^=�#��=�Qs�S떔��
]#�>U~"��o��P?�]��Ib=�������m�X6���pa~�c[`#��h�&�t4_����ؐ�#)>�C/>�,r�?��/�	24Kw��� �0�d��Ƞ�
��.�&�^ҕ�PY�(�����Md�%��%y�eލ3FM#9{������ub�ux�%�!����ӹ�0��_�T������A������ظQ�Ŝfm��jv?^���f�,�^X��I,~ej��:��f]0�l�����>��-�}螝�ǒ��V�f����`e����E�Z��ʢ�k�#���b��F?q����@x��j���Wc��,]�ćüۼ�>�d���`IWt5�Ftn�y2%���[0�_�}g��h�-r��V�F�8�e){2H����*��.j�9z؂~�K�̞�����rd]�oo�"��qNξ=ݑ��I�v��~c��p���?��I)��πW��������:1�����A��5�A����������yoC��UTk�".��x�X�uf>�;#[F�k�g�v �ԕ7�?���ɰ$��t�EJ�����R�R�0B�� D	�1�Fb��ݽь�{������������u]��,r�c�-to�r`�-�+��%K��������׆nC��[ ��3JKKw�^0�e�>8	����tIC��U.iI�)0w�W�y%as����L�#O�,�,��H)6��R�sϫR*�G��;Wcuԅ��u/,�E�ȴ����Y&�;}���I��_w
w��g}u{/t�c�I�Ȁ�(���>&|`x:h�.f��Y�~w����?"l�v�qMj���.�s���R=.��p��U� �Ŝ�r*�(����;�Hoz�9�O��z_FkT�*Ro4�ғ���"�����P%��D{�l�E�A��E��" =i(o��&�ZN<`}Z���Ģ�&�����\�L遆&œ�<GE%W�e����%V�t׷o��t�/	�N�H~z�*�=�c�;��#������MлW�5{��7�����4��d�"g�O��� �3�*�t�h�+����Xzϖ����1���37�U?Z!7���.Z\H�{x�-�d����Qū��/`0���isoo�L��&��aMq�E�`uN‏����Մ��H�5ت�ŹʞF�l�h���[	�NC�(�d��P�%�~��o�$��ݽ�z���6������}��ʸ�n�\Oi�1U�5��/D���Q}X�B��2d2�E�΅��0+��.����j�������ܥ���v���q����X�����Ǜ|$qM- �'q܇�s�ta�u�'2p�Wz#7�Le��RUh���]Y)�(D��v���c[.aI��w���}f��`�7�z3p	����0�g�oD�&�0?��[J*BI
��IL�Tz5y�qC.s�颤�_�R�y��.��%��W�am�Gv��ҵ���~c��X�&G���+�{Q���c���ez8�ˎ�^[��+���1�!ɪ��h����Î� j�G�g��su�n74x���ޭ�!����l��/3fbǇ���J�tc�#-����t{ܟU�#���ٿ$e�\#���mk����rǙgEz��qD��;�OOBW�쭣7X+��dUg9��f&%�SX_�A�`���8 ;�)K���ȁ�<Wuou}O��H�z�.
5�a;o�̳�����BĦ5^S&K��nv$��h\��3�2.�NZ띒�("d��U�_/Y�����8ռ=���8�,�L�kE��&������N����t��kGG��P�W�D<o<��s�Vrk�[1^{���w~���>'�]����C�벨5�o#+��Sb�]�8�MCzl��	��i�V�k�����'+���K������9��3������WP|�&��/�땝gr]���`�[;�$;gfԸ�_���`�lR��=�FG����d�5�|9��֑ˇ� �ѹL�(�����#^k�߀�L��|$se"A0�$��=c\C~�uuą��1��ٙS�Z�/�M����rs"?�K�h���%��I��s�I�S�%��B��<j��N�AIV�E�[z�����Z�������"�;B�	dweq�|w�D��9پ�ЋYX��ż%]�۬x�y)���ꢤƷJL7w��`��{Į��`�� �,�+Y4��YY�gZ�@�T��Zaa!n��~��O����T-����|xX�7���=b�;�ڥ�h�`#�Z*�m��(��`�����N���17p�m!��Q)�q�g� R�㯏,£�ƀ�φ.�!8N0U��	���^(�m��\'�?�P���]c�h�����?\�|B����	g��ͭ�Ƨ��G��b�Ճ�y�Mw�O���y=��0"N�̫��Hk=�~]ҩ������I�;t,�cҫ�M���JiB&��H;�̕����`�a���"y�ƣg#g�k��1}�

�W�7�;ӎ��Y�͕�~0 �;��Yd��&⻯p�R��5�pq0Ѕ#^			��IW���L%��{E��z}B�.<B���cPd"C����������sq�@�9� �?T淰��b����Vt�+>K i��ȧT^���?�*+�/s�ژ��L�e)Yb9�苣�aH���ȣ��|��Pa��s��颣�J�;:v�$���t�DDg0���j;z�L�p͵��p��[���33��
@��Ą^��A�&u�������I�<ݻ����{x�g���I5�B��e��$��Ջ�<�Q���6]iR��`NH��$�J�x�����$����xjtַW��d����|���g��*ǂ4H�5E�Ip�k���ja+��&�k�G��W��`�¿�9��c�ůCD�_@��)�@���m�/ӟ�ݙA�VW�����>fD�����	<��.i퇹-ގ�P�`0X��Lq��K�g�?��R�Q��ǝK����lY�+�R{5v�aL���GHr^>7iP��L)Gb	 .�C�1��="]���:(涓o�>�I~GT���HҶb<�"J����o�:吨�����eP4$*��D��$8��R�<R@^iy�55t8��྅����$	ô7���Y���5�޼y��+nxb"�����p!΃323[��:�+�����M)�<�n�	��v\��R<���^��OK���h���j�:��Vt&��nI�b9���s�ŝ�נ�$�N�i�ެ�<��^����.�}�j:I˾^'N����z/�q0vM��y�(ztgG���$�3��n.;��2�~�vI3��	���C���ԗ%	�W����.�}o���#'�fz9�0Ш��-�ƥ��h[��;k�L���q(z2��8Z�����(u�!@ѵ�`�čj�ێ�6.?�50��b��,��uu�JD���<&��}�=��ZP���mm/z�i�����O�3N�H�`�L�݁�����	 4А���>�䥆�a�m9-P�M�+�oo�#���ԯ�)�m9b$Z��hgq���]�&)��܍g��y�O*���%s"�6�2u�a[ �a�.ۏ�e�Ɉ�������7!��s�Dh��N{��?1�[�YK��ޙ��$]dX'\�U��>�t����ר}���&tf�S�<�{�|Ձi4�L�����j9Qa�x���bp���YJ#��[�28;u��ݩ�� j����ׇ]��eŅoޜ�p͆m]c�N�'ai1I[ާRcK��� �^�����0V�L�{IZ>�q:jq]W�q�}�����N]��>�q�]
��fQ��M)ymM����.�CW��xYK�{k��^,��Y��K�}��`�����QʂH�D�����x�e	�����Prֻ�qI" S.)��>9.�Uۍe�����2�\��>p�P~\z?P4 ���t���� ��u#3�9��7�prb�G��AZ�_������H�?�?�4f��Ru�"��f��Y���￞���%$K/'���3�N3�/P�]�{�s���涤')�q��x	^��c����'}Ώ i�m�N.�,��@��A�Z�Ό35�m�[�]H�$G�r�X�0���TyE�����#1^��z$�~�ߣZT�٘�O�����G��ЯJ	0�@;�K��dK����#�&�Y�M�F��.j7n�_��P�PI�
O}{m��h<	�>�n<u����
zg�@C0}���Ks�(z����ZѪ�.&�߷�4�����3]��hd�h�k?��@�{_���ge���(�Q~��`�ԗ:s�e�C���@�
�6�_��J�i��񙮁4�������M�<�B��Q���#�p@�Їyܔ
 �Ē3Jb����H�ƞ%�5<<<��"���Pk��8J�^mRz��0"e?�J$ć��$�MEM��LD^��V�lv)�f3��V��fj�K�#p�����i}�jG��.��t�=
D�
���K���������)sF&��ϳh��^���~q�	���3����q�}�p�@[�UPPPf����\������D���o200�ʔ-3�"'�������P���p>�%M///�7TUU}��0j���e��N'|ϡ��d��¿�[�1}���@��v	����o2�=ԕ$g�ţ����gᄑ�R;���o^{�$�v%��T�DJ���6�}h8����:��7�<��؈�8�v Pꅖ�FP��钮*E>�:ύ��k��8���~��pV�Wӵ��ܱ��S�Ò��ܚ����S_�p�|[��2��/�Y����G��{���y2kx��xb����)���iӢ�������L��4�͑ۖ�7�~h�l�"�///ŝ�_d��>q�	��]����jҙ��j[Z�#X��-w�T�ۀ�&��s��"{�Do���m�Je����JU������օ|%��/r����WC^;�.�J K(��+���%����Jl��)1��������_q|zKy�Z��'nó�jl2w|w��<�,���-ǋ�b���&� �}�u��}y���c#���<��av������� �.v���ϴ�~�W~q0S>���=����k'c��߿_c�D��`Z<�Ԙ5�#q?��\snn�n`	s��n`svrx|���G�D"u��%lmm���ɳb
׃xĪ�	��u����(%��=�5�H�7U͒��˃�rv:����4Kpp(�$�����	��A�@3յ����O��@`ӕn� ��w;/�d�O�v��B�N���"�@��>~��bꍓ�#K���]K�=�w�b��}~V�ꥡ���^&4�pt�殕�nx�a��OW��:ʯ�:�$��2������i��g�d�,�>�e�b}���;���̶iY�J�^�-�
oy�!���e>�ܫ�v�9߳<��$�`k�V�?8�w��s�,���џ�'l�Q����?[���s�����{yM�	jW��d��R� �'���f�.����_��W���Z�5�\��OZ�����L�,�{�\�$y>0z��+x�ɪ���v��������`��`Y������S�5�ĚKK�(��R��{�G���3�v�:��`��7وSb��e!w�Z�V���O�{�lư[�沣���+d5��t�����/8H4v��T�E�	�+����/<rv騛D��mq����$8������ۑ􂝋�C33�11�m{��S���Z-�%j���⚛5�_�{xT���<�Y4ܫC�(P� YH6c��{�~k�.�����`#"���w�x�zw&�**�lS�o &�Iy�[�?���%{]u�r�j7j����q���-��y�񍏖�������%�&o16��Ck}@^�O;3���>��/@q�$	iA;�k����������4�ާ q��n3T¦��ۋ��$S��b�K����̪W�TGB�2�v,��oz��-�S�.=�?������H0j������O��Ĭ��s�]�㝹�o�W�n�R�؄� ǈ�zp� ���Q.����3��E����rvB��/-�����M��)©Ԇ����}r�>�'8��t%GI@�2ܒ�V��CR���ٷ��A�+�6�"�(1@|����|�����O��� q�ж���iFpI���0(�9=�?�  ���!�j�`�,R^4��``b��?Qe�^ڙ�}������]�
��(���744�y��TUW;��R%x�O������d���PܒK�^RcP?��6��h�Dk���Vdb~�q��է6��6a�h��K(dٲP�x��A?����r�OS���(]_޸8�����K��DoT����l�E*���gu>�7Rڝ!�b��X����~�䄿tO>X3=����f)��v��ɹA��˙��=�t�b�c���[�c��D��D}m��V ;�r����iX�e�g؍���##�DXn,9������D���c7ww�Ǝ��[�����C��(z����/Y{�8�=m7��f�%��wܧ�@OϚvy_,貾���릲�J�RZ�{��W�KE/�뿲����G�P<etv��$��fb�V1}(���m�R �:�L	kF9[ x5�b��psE��0��.�ʍ1�ض1Qx��!�w���܋�����q/�-1�c���9{�"��������2�&qO)f�=��S�\�<�"��m��	B�pw��XYYu�l�V���t��j$��)��cr��~Lf�s��-ҕ7����K3�Þi�!h��RE�Q��H��l7:��-���Zk
_�/�����>�Ը���A������y#���Y=�}���1��B$��鄹�L��lI �'#`�ORMԍ�
J�a�ʂ���vn��vJ�F���$��J�K��/3n��֦!��J�ɣA��$�~g��㿍@y��<��Q�7�p�5!RL��7��X�Tp�׫�|�Q�n`��ϧ�[����Ɲ��P�����v�8��W9�T(3-����m\0�OT$����r�����K.'��$?����%8�����/��Tˤ��R8�-�4�9&���o�6��A{�U�S}���T��W�0�2��N����r�O�s�_���P����^!G�?�݈�t��iQ��,�Ey�
jx0�2\i�"F!���l���/]��`��#&-��`ebaA����'��q�yW���qW,�Z�Y GFn�-��Fσ��!�`���ũ����vv|	�z55O_}n7�Y�5ITΘٹ��,�y���@�l;ۧ7�o�h��l�Ȓh9�啙k��څ�q����7�7m:#Ѻ���3��Aj�H�����uC�b!'Atx}xQ���؎�]΅��eex�MG���`�38]�iv#"u�~㾔�4_�m�X���w��[���3'V�u�O��D�3�eƿ�9$sM4kx2 4F�\�>"�pF9�x�������<j��[Y��<�Fb'��Y�4�P�#����{�cc: ��a�Y�ō@2�����w	���Qs��xx��)4��aܠP���`܍'��^-f)F�9-�YI��2 ���!�s����A��98&^�j�v�3��T,�\�vy�f�[��o@��_�y�$�(��з�]k�rB���G�g�dսl�z�an��;���x�4� Z��Ms��x*�V|�썄W�/�ˌ[�5���<�{��%j�fP�?MG�v���N�bbGǗ���^p������PiR�--�)�>LKKK��c���N����)�� j�����wB}q~I�K8\R��`���9d}=#n��ή���`hr�g;9cn`� ���pD�� ��)�J�,u������S�V�Y�VR(~gu'���W%���@K��$�y����M*�?W"�g�+�*�\"6^�Y��{.m���ʟ���fLN��b<*���o��d~M�3�p�9�����o�]��L��]p=|��K�ϴ*N�~϶�<Y���7~�$�:�~V�R?;?�j`Pbrx}!�E�&��oT��s�1���0������UT/��N�x������ַ����Xs''ʶ�6V֎�Aʐ��<EvI(555�G
4�������H���4�'aU
�RK �����ݖ���=�}�N4ų~��Na6�q#v1�v�[�zҜ�u�����S�')XR����z���r��3ukx8Ť�o(��Փ8Y#zH�ɝ��wz p.���[�1��B~+A���A�Y��3����zw㿽5H�,���������cL��fmW+�{VP�8Vvv�BQ=N5O���\��֖��߿I�ɭ��4�]]��{{�m����o��wW�_;N�7���������L��C��agg^O�<� �ITT��h[;;܏FGG�lRG�g6}e��I[t�=���S��u��|�� �A<|�4&`�nM~^>�Nà)�v�/j��04u��\:!�t����Wo�6���9����!xyZW@7���֍���b��RC�&ҹ�V4���3av�� ��s/��1~���Pwd"RT�_�u�Ay�q_���,Z�����rb�9�R����w~���n���X�	uf'��f��.��/��U�����l��{�����}a`g�g���5��͍&;;����p	?y��9a�|�㮤��p>|4!�XvNNμTMUUFv���������I�0k����W�2{Bb���5�C�w��\�C����Ip#�dP�)��������27��I���Q����i8a���%�,�Ʃ�dt���B��`|{o����ob9��>����Ǔj�I*��A�M�J��� ��Y��Z�}�j�2�_�6A�w�5/A�Z��.�`����������{��k� |��1�������T����x.�e���=3�}�n�ck������^����6�mn���S� ��/3\�q�>L[v�ل61���5��ÏO���y��B����&I4����o�����Mݐs�M�`�_�:�B��~����eT�;^�%W�}-x���0������L~�N���rCc���L���b�.Z���^��b��M?j�L}�M� }l�p����F	�c���)�|��H�Ph�8Qm���	��{��g�R���L7�O���̓;u�� ����[  �����(���v��	���\�4I����V��%t[�z�Rzy�൜��ȝp ���L}|� �V��)�231��T����K�|O��n����2X�gb�R�hV��*�1ڦЃ���TZ[k��ϖ�f���b].�Y��$���I�D���'�4%r��:OF�����GY�UR�����(7��#Z���xCf�[i2�D�^!Dhy]祊2�q�@R�0���ev��v�M��x�� "4ѧ_�wc߽�"XV��Q>�9؉Vg�Y��K�r��օȿ=�+䙠n��3���h�g z<"����-Ƈ��ڰ)�*�1b��{�6bNuk2h�ޥĜ��1�I.�.@�2[�/�17�eB���S"Ω�Z�n�;�H�آ+����W��X�U��eF����+.Z�*ff��6̍T�ۅ�$�)��cܑS{��r�i�;)��y�3�Ky����BwG�����#�i�2�Cp�i� ^�\oU�r�q(�K3E{�n�?�����"�G#s��.
�g��;�
�� S�h�mV��5�ev/v�)�eP����hR���ڃ��Q��-��gRN���G��M8��Y/qGrWGYڋ����Q���iVaֱ4����^C2ˎ��A�*��"�Ww�2��-up����,L�u0+!!x�z��B��-z�^o�*4�r�R'�9o����D�g�怯�*�}�i&��[�ۄ�\�o��������3�z	ѭ_U�M�Tl���Op��F��^Z�����LU�u�5\��_,H\,St\2�d��t8�Y!�<���3����/�������~<�?���D^�Er�d0�C�h���}��o86-_SJ(W3�0������z2�f�
�R�L��c�� KjJ�w�C�EWz^g��-K�t`k���X�N�����d G����}��"��ڦT ��?]��#�+s]��Ƥ8L��#6
��'��p{)�ݎ�j�v�]��b
3)�V�O6G���O��ud8�<���gb���fa)kM���R;�mq����-�Q8�Ӕc�>d���f��a�(�I�Zv�c�^�<`���큺�W��N�Y�2Vo#��V���뭊�3��
=	?�O����a���:ϢP��y�E�.Õ�8t�>�;��1�{�-k����-6�cAq����򞎕m�*����l��Z�Ɯf�Ŷ��!x݃G�UA(��;n�"AC�����Ût��u�"3%İ�����/�'+��j[^���&��%�]��4�����^Dl�r~Uo�r�-d��)Q�����bgI��I�1�چq�g�i/���E+nK��W_ �@ɢ�̴�z� Y�}��	��n(��=��E�%rn4L�������Փ��f�.�0�G_�8���?��O>}~1Fr9v���~��A<w#=�<�l̲�݂
�9�ŐQ�a	�tzAE�x�6G�u7L	�<��o�4N�z�9k�� �Bf+k� uիUk��z�Ս��瘸��׫eKH̦?��Y>�O��c�/BpGŠIak�w>)������8b��Χ�?��ç��� ���6	a��;4YZ���ְ�ٴ������}n��EpT��R����8(u�
���<���,��Z��`����Tʇ���9��nJ��I�C>��x.�{�*�,��8�W��X$��ίmV�#Pv��c�C��z\M�5�@f�{��\ʓdr.r?�%�U��#O�����-�6�OzRT]�&�-�i�+��O�(w���vA��z�K����[����碌��I�'�Y��Fr�-�W��[1ϳ�SM�GjȦ<��̈́s�A�"�l
4K�1���S�֒�fFj[�+l���I��R��Ty6���{e��|��3�e3��-��T%�������7<3��Ŗ&o�������>'2;���
ӱ��n#Kg*���3*�kv6��E�RyWy)G]�Rj6K�Fސxh?0���?{�JҰ%�`r|�2~�lNX��G�Z��$R�i���g��ih�0d�ȓ���IOy���0M�q�F�����eȆ\&� {ɗ�ٷ�j#��p6���0w�Mn�#�z�&!�:����,
�G�;�T��_� X��i�톇QϚ�.�@p� �8|���,�Z�v=���C�St]��. ݀]�|7F(�ܣ<�2�/ ���2���w���6�Q�܉{��Ơ��g�=ρe�<d�f�,�Na�.�\J\��4�s�|I&p2��]_EQC���1E�*�����]��EIt���I�QB���i�M�O#��eRj���}
s��>���Z;DJ���0K�(K�E�L��O���\��7�`��\��
I���8�E�=0��	G�w��|kQ����i�y���ʗ
h(��h��İ[�N�@�t	�/XH��.�����h��g�z�`��U��u�$��T�q��3BK��#g�I�`��ƩǂV�)�!q@��ئ���kN��=N�x}�sr)r��K+!���&[/�p�?��6�D�)с�,�M�f�͍U%�( �`�E���+:����`4���B���������%�zUʷW�i��in��D#)N��x�h#�uFk����x8��*ulIg���/�?���� _$�L���w�d�8����S��f&F>'�|>��ǃ;$���?��N&�
drS��~,�i�٩4j�i��o(�������	��*���/�FR����k��0��-Q\Z9+�2��q����!��3];ǵ���pD��U
�7��3�T���E�����X��|��V�W����3����{�H��-�+��tڑ�EfhB���1�D�eW�ƭ'e=gH�qI�?4���>}�}>�n�Uƛ�[�����e����]��/�M�~�����fu��׾h���Y�a���jՇ O��<f�<( X�`�zs��8N!D�,�]��>c���c�����#�b�I!�(��~�C��Q��������$<dUgV�|Wʓ�qH�%��u��GX���}�ϲP�Y�>Gꃝ8����g�4�z_L뼲H���^�x�7`V�o�*Q�!�ؘB/���8 -�nXq�Eg���c�ok/�nSu2ɸ���QC��Ee����&t�&���T%;���>8$�@gAV�=o�Gj��L��g4R*(���=���Q��k��s���u����+�<WǷ캢�袿u��:/��w�A�Ѿw&���s��nCL��޷��L�m���*��P�l�^�����(�)���%����ͬ��e9LT�4ʇpH�}x�'O�u}�e�I��S��Sy�HO��d ߬,���븡j)�}�-&�V7.(�'\�x�N�>٢{8t������k��u�>��X����La�y�RZ��TQ:�A����լ��b�l�r������Ѥҵ��I-���@���K� tAAE������'��M�@ �T��ؚt�R{�9Lk���U8�j��E6G�ף�S�Ҙsa|��C���D���P{��򩓬A�-g�-'���=u�a���}�%y�XϢC��,��s)	d&ݝ\fwYD��c�a2=��Œ#x��%�c<����g����no��ӮE����;ʻ�78���W �Y��a��}�yZ���.Y�^��7A�B�HٱST+�A�QT�1v��{��
��f_�t�Y�M�P�������.S��	yF��D�LH���޷C=��\��:��0M@�f�]ǌ�XD�p��O�@B�I7�r��<u$u��[ʾ���=�>�K���)'w<�#���6�^�cΟ��������Z��?	���F��
�&l�J�ަ��<o��i�aW�Y$�a�Iԍ�%���W[wI�;��j�D��e��V�o�o��C�7+��/��R=�~P)�����^�Za�{����KE�QY�~���l%R�P�H]X�W|�88 �4K�}{}JF�Pʭ�����p}��-6�pm�[s|�e��*j�4"��� �Ir��Ii���	9�)׈�y�M`B.��gq�z&�{����f�;uP�8�=-��"W%�}I��ӛ��s��p!�hST��5�M��Y�w�3�f9D�%�z���{<������'}Hf��|Bغ��=>��R�MN��ǡ�y2�#���+�A� k�	߄`T�)��ל�?���Gi��2\b�^��{l.�S�W{�y���ԑ�Ng��Tz+�,������ץ�Iн3/Rxޠ�q�A����=�����[֕%
|\��ꤝ&N�	7�ڦ�X2�u�o+��U�/�re5����n�i-���v=<�-��j@�Z��$�&�W�4B)�����MtȹG;�e�1���3Zyo��#��$�>�^���<v~pj�&�����_�f
�**�����6�ŭ�W��lF��^<�[z�~�xU��\�c�8=��hz������͒~�p�����&�����7�]�i��zA�l��7S�`g�U��k��,���J�Z��w�	�E[I�|M��[���S
�2WiWg�d5�Z��P���۪���[Sz*�U��l�Sޣ5�$����9P����+��,�2�}�;|���wb�AdIш��S,�m��w��N��-���\���ue<���+w�I�Q{Q�%+]W���A��Qe�w�}�@�8zv=�qjG}���w��V;j���(屖uQ)������������~�"s�ș1�6���"2�Q�{�z�$�[x�I���Gg�3�����+(�l�9i���'�s���xNɎ%�3 }��{�Ǘ�RҬ��5]W�����Yz��Ӽ�q9�=����^"JwE�-�(k�%M��#in��O��!q����q�G_��E7�CXJ��6�f��ϳ�F������vG�L�wţ��Wo�xwPՈu����G�6��p������;y�*��O׽
E!�y fl��و8cN��������N�F�����>}i�WR�JZ��@4��`��xp�C==�`u��g��E�U�Q��N�|�ƅ3ޫ�xl�+`c����x8S/�UEc��9.����� ��H�fg��L�z�!��bh.kBݡQ�/⎣{����;�L<Dm.\�X�XP�#KIZz&| ���9:c����A���&G훫�2^,+X��]f���E���ހξ�N��<Ҷ���^�
�����V_��%�<��^R� 5$�,�O&D>�m�st���Y�%�`t��W�S�P{�cC�|^�Ig���k���?8
���~z�`)���J��W��R ��^l�<����)�5c����M�;fN���/�ܧ"Dw[-�?r@/*|�It@�~G��T_��v�J�4�瞗3c|�1J4�NS�[N��W��hz���_jӱ�u?�rIe���^�6�k��o�9=��j�r�ķSK64ǉS�(P�cu�Q$Z�%ŽTmR鴢2f��K9��?�!��!A���|3Su�dō�w�7�~��oz+��~y�{H�t�<+��C�����-���q$k5�O������][ge���R�Bk|#����
�:IN�쭣��ma�{��!�~VN�Th�~%-0�ƹƴ^7/c��<o�`S+��L@��W�O�P����f1r@4jI��M��E�˸\���7F\��g�s�0%��!n�piK:!�@<�*W�:�2ڲV��Z�Dh�h�G��EhV�m险�?����%������7���CG�|
�j�A,�>���yp����S�p�����.���ڌ��Bi>��C,[����F\z�n$����
W�yD�bIhz�uӵ�ۼ��w{BA	��>׻��� s��5��c����O{��L��b�ڹ w�HRs뇹{�>��1�]'A̛��O��>��=2G]o��]naO��J�ٯ�[��&��pyd���) �.~���.����s��w�˺��e"u�7JRd���������t(;���%��zc��Vn�qd;���p}���$���#M���|)9D���|�u>ҋ���$�ն�)���<i�x�_��-/�R��Y������j�_��>�g�%�u츊a��V�uUg5�hSXDZ�"��̤�����xM@;®�d��\t=���VZ6���b��9��N��/��U/GІ���#W@~��U��z+�2Z���3c��w����`�X�@q?)Y�9%*{�hY��v��+q��>��o�3�ܢR����FW��b�!#�.���꥛�*�>G+�n�~���zf����S"�Ց��ZӛnMu�2�K{���d������0��eS�JOQ��U��e����JG�|B��d�����8�ki#�V��P��/�b�y'�HX
�vq�����������?4�W87�Aj{��'��d�w��ô�;!E'���i�)nЧ�x����m��I��%��s�NR�JV5��!�����ԙ�U3�ɹ[����[�XK��I�h}�@����%��}�6�sz�_�Lc����O;�-�(�.X;�8����9x�z9�ؚ,�2�ݿ�(��ޓ�B������4����P!oE�9�\ٰ��ii�d�������!x����Y�h5C	$b���Ч���8�&��b�p�4/�h/\҃VumNR��IU�K�\.m%�V�����1'��D��I#췜qW�ʵ�j5��/�w��'0k5��E��8zd�Oa��x� ۍg?�yI�"y�u�,���O~VV����`R�,��l��f�f�mo@���"�����l�p���_�|D�[R�4�ɨ��� |Ơ[% ��C�>GP�@=ݖ4�}�n�U_Hq���,��/�e.t�������:D�����d�$�Ąe�q�������[\����}�����k���2Jo�Df�J�ٯ���u\�=�<�����:��:n]�.88ː�8%��M�1�p��(��ϊ�Ua����=ü>����l�J4�i�7�&}�>h2}/����� ����fbd�e���ܡ��r�MHV�[>����[X'D��%��^�e���{��.U�>e��?Dy�p"�2
�B��� d�Fz,���.�TY�<ϸ;�DC���GW_J�čc�>H�Y$�$с�r
{���*P�QA�p���3���L���)����#���g�S,�y�4L�H��&7lO��HV�ũ*q����� �*&6"��$C_��R#�=nHY�}%����uB8�v� �@u������?�tB����ѺAs��f�+��^�HWj�3֏}�r�Q�E+�Dt�p8.s��q�@�c����8���x4�4qwZZ�K������)O�u~��)uL���F������� �]ze�K6���?����lw���e`�V����Њі��t�F�iq�"�_h+����:&��/��j�`ῐ����?I�P)�Պ0^�Rv�� n3X�r��o�ny�!&z��|����M�*�|��m��V�[�q#��|� 1��#���Xc���ms!��h�<>�* �:C^�)S����x7x����/t�KA!��	�(.6���i���ރF�9���ϳ�O���gL7��}�"u�'�[Ѝ�Lb�E�[�k64��?���O�j#����roX��$��o�M�㱯�w��r�H���T%p}bD�VO een������O/Y&�nr��?뎸�D��΅0�{�o�㰬_	U�Ǖ�p�ӄ�R����w�{A�ܶ��)E���jE��j�����x�ӒR�K��6��3p��*��̫�e:��\�[��3��T�bz����[�%����C|íO
�Qϐ�����b0����\2���(Y���<#>�V�8Y$��X��E����N�`�� fy�4u�x�<*��y� �!H�2�ϧ�'�W�����C�N]v)DԮg�ٙ�ѧrSN�QlfI\�"Hy�<�|��G�;����	����ra�-\�����J�S�Zw��;���-��m,xZt�`�3�ɴcJ��]��5lF=(������ʧT�R��������;�ex�
�"GO�Ai֬^�R����R���	�90�и����4���Ad#�P�Km�~ �JfXF��!)(<Uhg��P�L�ڍ�Q�kWŇ���[���N.�v3��\`.Ckn��R�������5C
>߹:0��wT����ϻ�0@�q5���~w���0O�d5��埅��ֺ%���9_���{@8g-O,1nS>sR�>��Ѕ�Ee �P���23}�:�|)��1�нO��h��Y�m}�I�l�`��
��E�Te��~�g�W����ꭣ���7P�iAT�Ni�����n$�A����CAJi�a�B������]��yך�X�����~�}�9�,_|�;vȔ]�ؽ��G�&�t�v��f�V���3^�����v,�r�xo=�-�i��һ��n?���B���B�H����@;�ү.�T�>�O��Ɇ�9�n�K�2f�$W+�*�>�	�fQ\=��R'�(�M�\I��η���v�h�<��Ag0+Zs֔hCXw�1b�?�@n�{�vv� <�y<i��ѺN�"+�!v��r�!���lk�p@��7�Q���E�k�=��ƿ��L@�H3ߌМO��FwH���^R��CN�#nn"�%wt�=����o@�-����}�k[�o5>�<���?|^^��H|��ap+�!K��2m҆�y�d�~M�Ē��+Ih�.d&��<��7���+�c�b���?G��]�
.���:��u�3�s�K3��q�dd$4]I���ϋo^=듹��}Hf�Y���?���H_ϗI"j�����`@Tc��񈅘3�M$�m�1��=���! �a@�u	f{��G�]�
R���}96���i���sQ B(���\�߈�LC��w0�7�u
 i�V��\�+�8mw:���揣�|�Ԟ��bXh!���k�=V�O�9���V��k�v�e����-�I���(Y��>6���,A���F^�����C��!���R�����'���'#�W�"+�ْ���b\�}$��d������VH���~S�b����iFş�4�h��Ӗd٣�69���.�gu��Z��D�ц��,�=�jrw��.��]cL��u4eY.�[�D4���K�+8`��wI����4ŉ�Y^�.�s���$
�K��o��}û�=?	a����50����"�
���$�!�����f��K�l�?�IВMm��F
��?���4�t��Z�-�d��.lP��{�ȖT4dg��{y�3������v�����o����R`�L&�˗R����/u$fj��-����Jɯ[�u�7�i� ����g��͡7Gh��.l��A�������߲�����Y#���S����(�����`d�-[�j�Nڑ�t'.��Vҹ������)qj�����pw1+�3���z�	΅��Byl��~���3\%qEw}��G���(���,Um-r>��BH��P&d�2����@�����8]��J����S���lw�/ڎ��H`�˳�^F���׆����������}�7j.�R�H���a����L	�vr�k��Jf��EJ�̱LŲMN�rjcz���)���. [��d���^R�K5�6ms��W�Mڴ����D��~�jmB7��(kBA��?�K`��a3�o� ��bC�L;���ܒ`�t��E����0�]D�n��}�{4� 7�#�a��ɩ%�T�!��!5�Pk�1"���)h����C�pZ^�Ʌ��p���d�OV'n��5ǋ�xOM^秵&��&���u�����X@�u�sg�>M�A`u������&�X]7�������I��r��U(�y����8-9�Qf�4<��-4�V�=��L)�%�]�xQw�H���i>�I��y�Ö%�$�W�u� ����`���
�����8y�{Q���҃U��<�̘;��sꁟG�tZѿ�����O��;6�0ި� !�;�wH�<�m4��.֬��nˣכ2~Jg`Y��@�ö
Kx���ϕ@�W:-�9U�{�1���_V�:��^КA?�j�=��$�/�1n��K��3oAZ*�QX�\�������/���J�����}��t
p*O�&�ҩ'���!0���H�ےc+8�NI�����;V�ms(F�S�r�R
h�m�zR�!H���~��ZJO���>�� �ݺ��Gǵ"��lgK�H~(������(���x�Gw��A����!�1J�sD��3j��IҬ߬�Q���U���r8O��z�^�{XR���Z���Zh��0��{�#�e����P�6o'	}�;�`/��j�yL�I	Y]�Ә�h0z�)�I�E�������x䤪�E�c�14!ݣ���n�p���(qU��9�56�t����"� A�w�������}iԢ-e�-���?2F����!^ǟ,�4U��j�l�M����^�S���V&:�V�D�����a����5H��~��v�H�LG,��>$?��,5e'�t2�N�/�m��@[����:��lk\lc�d�-��N�^����� [�<��Tv�w�g����Q��$�?�i��'J�0|����P&E������j.Y6��J�����^�J��Si�2���+� Ф�'��D|��ܹ��z���úN_ƛz���j�>A6x?��8��nxӺ���vH]� �Zv{����/�&�b���a���D-�3]#���xa��x(�3�X3`��Y����n(�$]8��;!Oֻk&G�)?yx�c=܎���?�C���wY������ag#�,��xz�M��&�QW?��%��6�J�]���w�\��(��`zu���{��y������Z�8�c����-R�Ӕ���ݔ��z����:�F�!g��!D`��&�!�(Ύ�F�#u|�; ��	�/VT	N�g��4&����Q��(ѕx�'2�3z�#ch�Q�䵼��J{
���w�mA Lg���I����J#��L�c�o���#�׾,k�Y�źq�{2�Ɂ�����z���>e��</ol�{� ��eq�t�|<��Un���T�Πz�*�ek�4��roa�mj9�\p�c]����2�W5Y�m���Dw�d���$|9g��]���/w��>�?�Ń�	]�V}�+�D���Ÿa���6���:�1Hl��'�h��@��3]c/eY�_���5��k���V$�(lA]��O/1-�����-�����b �<�����3��X5�:�:k�3ep�%5���}�ɿCn�S�;&9�ߡ��2�O��oi�6�����t����Gfp��.�[�gAa��s��������"o���_���F�<�>�gU�J�v"j����
,��d�*�R8=��k�6����g
N�^|���[�5&i�b=���z=���ƣ����X�$�	���_��Ҟ��I�~b�W�{p5�lK�ys"aruP�!?����l7&)6Ң����)"�=�7��47�~����\�����"��ގm����ZC7�ϖ�׿Nc�3�!7ߙ��e���9%U^_��ɊȄ�<ޔP�+�֟�o��S�g%I������3Z���GT(~�I}��?N�ؕ�R�?̚��栫ߨfwJ���Nt-����{�J{E1PCot&^���$��o�b1Y�n1������wx����==��X^��7O
«��9�b��6��V��}�n[z>Ps�`�Փ��l2P��J��
�J{n��@��q���ܛ�F��F�P��H���
~ .,�)�s���j1��n3�d�J1˖�*�匏m2�;b�f��V󟗺����h�������ˮ��
@�3���Y�dJ�$����t#DD��OmO�b��X�j��~�r.o#*�	giz7D\ra�������:�����������Z�F:U��ʊ���M�|�Ws���:�!w.g�Z�ۺ�
�1�)Sx���a��?h5F^ D���7�X]P��#)h������i�1^I0�$$4�dY��k�vp�>�Y�FLy��] j���W���>��=)y�q~GSL'�Gmqvt�st��"�C�����C���`	?�i6,�I��󛲪���A)C�I�>�
����eFW���i/̜=,�)�����fݬ��쾮�fP��F��b��#�^X��;=�M\������`2x�[�$���4�{#5A����������2�.I����2U=5�Ͽ����e�:� Q�ok'm=��n�_Z���pj�1 a�:U%}�Щ*�I��5�~UvD�5��|�'��G�
���OLrf���=�.����ZJP#X���b��Zyu ������{z��>	ʃ��ոG?L�G-Z�H)��i����AS�Ύ�d��C�G��dU�}�1B�|<��	N�+X#�&㉤��}K�� �\گ�_2��w��]~v��3��q��ӳ'k��yT�'[W[O�:r}7�� e�u�2y��/�.�l
@������.a}�]���Ao���n�4d�S;��*�4̝���>@pN���y`	���5r�O*����t�{y� hI��?i����$���D����n\`��=�2+��/g�^��n\aoi;~�_��Fd��^�	�G���ꄰ�p��Ə1ׁ����9r&��̺_1 Cﲢ��
&v�L(	@L.���%W�13���w>ZO���9��(DK���"7&�i@���ܿNys�fj�w ��(��g�rnd�R����8��:��������>�J ��Zh���h�Di��ӊ=T�7J�{��.�(jV�K$��!���`��������3"�.o�"~����ڤI���vlN���|�0Gz���R��:���w��00���@'�,���!g��ى�-�TI?�l�����s���O��0�:�F�����Ze���_+�q�K���WM,ڮ\�5�ׁ0:yå0���Vͳ�%��Gã��$qJ��x��]?��I� �^�_�+pt
!d�ͱH<����	�W{�3iRS�/uq���F��u���%��(SNJ
gB��-N���y+�}f}�zM�Pm�6S��n( �Ϣ���+�i*��g7�� U��d��(���/�=5� �WJ���kp5����K,I�+�׈s=?]�Ճ�z�q��qbF?���;��3)YpEk�p3B��ތMR{�:��d3�x�,?�����s�@���Z�aw�mwh=ȡ���!���V)���`Zntt-��Ώ5�fw>������o���4lm..6bBjQ��ܔa�9rt@�x�d��ۋ[wlOY3�l���5���7�
���h�Ǉ7�p�������r��?͹O]H8VO���vb����W-��L:�*�oT���0�,��W��ߘE,{5FF����<e#j���P��>�5.U-�������g����1���@�{ZMp���f\��d4٧���y>�J1/I_P�D�1z�����m�~j�H"N3�q�t>Q��ѕ��5b,Dkʄxy�ɓ���똌�#�ǡ���t��"�(�~տ:mxE�MH7��=����Qt��ѝ=͆2nD��QKɆ=�1�UKör�'��qJ���
8�Si����*t$o�s��:�~�֥N�S��4d�p�xD�A�|�}�W����W������':�E���FA	��o݅v����{~�K���z��#�(]�J��x�t��	e�P��~�B��BP��Y�9Hj7V��x6*g'���\����>�U�}��5����_���<v��סZs�ڂ�T)+L�AM�~PH��/�����u։�j��y�?��Pb�=0 �L ��G���k�������TsR�t�p��X0a'�}��4I��T�|ND<i�7��Fo��������|7�S�y��?)�$�mk��R�L��Z��)���z/S�o����8'X��G�6'�SQ2Ň�iy�ks�S��&���Ƌ�߈|�v�3��{p�x2�,Z�/s�8����b�Z�9!��\N��������:{�s���~��⹘6���2��&N�{T�Ē	��hV"�W�}���r�HV9Z�$�*��yֿ���� �Q�j��I{���z\��%H�Wx-�7�wLKV���4��8bQ�j�L�<J1rq�o��<�d�\_¥������i@�����#2���"��Jj���]a�%���ցB�Bȍ��K�E�%�/3�a��E���뎌�ж�ݻ/G�m.�yA����?� щFD%�]Z"�mda���P���"*$`<�� �;�9m|In;�1�{�5�&F�Ys�M[8��x¸���ސ�1��}z���s2ȶ)jcfQ:"�=�]~[��!��];���d������?��l��.�����*���H����a�����ݸ"����<�,��s��V�\���oO(�=¹��,)��J} q�2o�����>9�)�|BA^����cjW�xC(�æNAa_���md �_ZS�����|�j���d�|�(�=��6M��!_W�o��ۜ�a��@՞�׋�෠�bv�`�Q��_--#K���9\dt�j/U;j�Z3F���]�����o_E���A[�FQz=�&��[r.7�9�\kG
�A������:X�`��~����8�g� J qx���X�J�nb�_*0aU�m��3?_I����,s�I5ͼV�z;����^��3)�x��s�V��K� �Z��?I���.!b;���+�k�R"�w�jċ����	��I'L�)5ZT�0�F��=�Fy�����o'���������� �(SB���D�##�;T}��v~���P���̹��/�������U���&�J�^�ނ��?� �.q�Ʈ���>�)G[�ϻ����LGke���q����\�ӍSϔ#X�1�U�Xr�1�Fɱ�:`\nx_Va�b�̇��􊻲~��i�����!��(%>���o3#X��ʙ)���jז�����߄�[�wtg9U�}����.w'ؘ]����27w��(5�w�缀_7�U��O���h��a��m#���ϕ��̖qjG@��a�,����#���>���A�v�BO@L�dV�sl��º��q!��z�wI}����3l#$G,�8�{,�����o@8c3��A�?�����[�[�m�_n\�oJ�7�S�>��[�N=�!氏��iq��Z�%a�Vh�����&d�^�P�[��HF�%�f�cV��2��E�N���c��V6p/������l�a���[�/��a����������[	2�ka��k��f��;�j<s�E�}G�k�"sj�C��#��q�L7Ă���Ѱ���o��� ~QdC;L��w�f󏆍@ ���1r?r:AH�rCa�C;8�%�'�h�L�L����{*��o�@Dt�Ies���l�:�}�9�"�$h��t�NwRXZI���$�cv��ч����I�5͍��s9�B�~��m������O���I�Z&ݢ��v�U�Շm���[A	�0ha�8@���t��r�4�!6)g�L���bNyA�֝�/�s��^��ү|O�� ��L��*=�4t|��j* ���RxN*uŒ���}Q���봞*� ���v���mZ����v��ݦrM���U��f�1�����X'}��V��Eh��8Z��d��Q�Cf !���G�4��߷�`� ��R�{R=�FVv~7����|0Y��gEU���H$"ǡd�,��Cק(�74�b�듇+���>&7�IZ�MvZ��ڣ����������!�F�I'm�2Sﻡ��&�w�g�kL�I�����%X���װ �h~d�s�����H�מO�7*�a�?���YV�rw��8�����7i�s6�E �j��4���8fh)��Οz��׳s�p[����\�u�Pa;-���X	ZX�6	<�*C����H���U�	����-a+�A��H�@ta�E�n�ud ��z�=D]+�u���^<b�%��n�
\t�_ܛ�@�f����:���O�[9������-�m���su�B�TO .E:)�OIP+�G$S�����`/m-�I�r��'v͈��ڍ��� ��D]�Y�D� �Z�v��_P݀Y�cCr��g_�&�#L�8��'�>��A��oL?"gE�ť6q�N���9C����e�����ц?)���.���S�"��96f���;[vA�/�IF�����D8e-w��9���:����O~��ۋRL~g#��XO
0���i�y�RW��	�hV�ӭ
�:���{���}L����`��4�HI-ڭ�1[��օT�l�J�#�2�X�v�#��z���`B�6����D-���!Hi��ɧo�f1_r`�����U@j&M�YZ�nٳ
�'�3#
[���p��8E��bT�o��f��ƌJ����c}��O�Z�b�T��HK��E�8�N��ZA�&cu 2 ���FL6v)_GF$-�� ~D�8߿��~j���Ů>d�9����⮡8S<��3w�~=SK�	�.���Oe���X����oĽAb	H��x�J��;�N������)�ݢL��u�_d_�*x�(ĝ~�f���J�Ƚj^�N�,��Ci�o����S�#�f9UX�e<2�����`�طIe��.���x�x�<��L�iz��;�C7�g�ZN�Yo�0J�Ț�P���*Y���I�>:���ju���M����t�������|��)&�w:L1{.?����׃���J���S�_�j���il��c,�I)	��Ӝ@n'?Q�6��(�N�g��ACw�M�ly?�3wûQ�fT\�����h��T��O"y]�"��⫷�=�m�I��`�1e��m�oh�7�W��*�`���a�?��>��{Ya�6x�msSz̵V$�'�u?�;����w(�
(�hν�[s鶒D0pk>�2�j�[13�E�%1�qN�zU��Z5����U �)�Jg�K̳@�An��`�ޖ�:p~eX_Y�Q5��_�y���>kEn���&n!\�]��l���G�xU$��3*	����5��!��~U����q],B��n�釘�4�n����Jy�ދ�W��i�i�{%���J�[�,)0���Vꨇ��8�bi��8�JZj�O��&:��z��;��Y�)=΢�z8�\��f7��������\���'��I}�'�Ļ1����P`�7QL%v_�@{��{� -`N�G�0���}rϽ^4���q^9%M��]�q��ܓ�XHmPI����[�(�[�L�<���^�䮊ܓK�)�<�]-K]�߻Or%D1�')����:����;\�4���eS����`f/Zvx�B��N�����1!��B�5>���_�y��o~�\����^�.�SQ�JFT�M�#Cd�6����I�T���%N{S�A�4��C��rX+"@M���q�{'s�Dw_,n*`�?��-X���8�ͻ0�e��ۈ�ܖŉS��Kqq�8�j��l���
�à<�F�ԙ���pE�NP��I\�Waקt]��4��+��R��I4�勆.�����hN�8�~����Ĺ��I�4l���x���Z|��/��@#�W�q+�&U+t\�Y���� n�K5��jՐ�6gS��0�N�]"Џ�hգ��!vU;����i�*�0�9�c-�	��\�S�W��%�p�?�z,�8��Ҭ����W+���P<I��ȕ 4�,d�_�5 k��-Ε�i�@0��	"�OT�*[Si䜁G���j�	���%�AE-��Em���E��"O?hB��Q�.�虜v�` h�)~�ôፂ+�#
T�h�`eڭ��CV�h��C��,��,�����׬R���7d��%��?��q-�>�u����$��<)��G�;�8���H:�c/>,�+�減F�KUf�D�3�\q�_5�p,��/̕KL��zQ":�$�9�
ޖ��v��� ��tP��Pc���6	 ��>�k��C��2nj���N��T���B�=R,ع��r�*mRyk���q������¡�~�D�pt������c��f�k�Ϙr�/f�ݼ1qiH���6Y�sR��p�Y��R��i�k�[�֦��x)jS���"��A��DD�*�F(&ob\mW��ơ��e�3��"GkM�m�ŸMc���ڎA�Xn�˜�b�T����I��CF$$��9�q=O;�ݘ�I�4q�\����*�7v�Lb����)�N㵅$o ����� �NU�'��D���3Ȇf%
��Z4<��FȣL�n�R�J�mG��O�:��h]�5�y����ۦ�Ӡ�����^j?R9��ۍ@Gɦ�U[N@��Z��W��P\qY����O)~�FnJS��R��P��^�LƄBC�l��GSN��9b�(��=t��DJ$\7ǥ��y�����7���Uva0�vc��Ѻ�W�ō|���@2���Xe�h2�:ǄBbd��%ic�tZWZ��J
���ƛ�~mM)K^<��_N�jζ�_gn?y�,�$�.��dW/^�1�݉ީB��l�;���k�`٪
+���>9����O"�G�0&�5I���Gm�t4���l��"��v4��_����'T8���":�v�C��O�B�R���L6o�c��r�z�ދ��S,��'�}Wҏ'��Q�g��{I���b��t �k|�u�AS��|�_݆��_��6x�g���$����[_�kG[���i��Gw�1��\��J��K�<��*�S������R�N����z�Q��)LE���(T��~�$����G�
K�lN8����=_���|�"���ϬW���9E���2���|4Ԭ�9��ؙ~�OK�*K��F�B�D�("���T�iI#��?U�	�ԛ��w���̽]_��t`�x��^c`I�g��IK)E�L���
qA�)���]��\-�ϕ��g�Z։�\r�PM��Y7�Y�C,B���� 9	:�dϦ����9b��z��D��B2�_ўK�ܥ���D��	9�]��|h`/�}�{����T�={�9-<���%����X̽��1����|�ʅ���y޽ir�.� �цh�=�+�ɲ��^%@E���r���a�zs�wT�����͖f�;����}��c���XFt(F;p�$'`������Q���Nbt��#���Z��ױ�􎀝�\��Tk���}��'U�c	:G0W1��Z��W_ �QCU���S��E��o�#*Tæ��9�ϫv���R�ߛ�?�.����
Xǒ����-N�Q����P����\�	�r�`H�:T�v��R��'%F�iX��⽿����0}�ӗkH�#�$����4��?����͉�CF��;F];�~'��_�Zo)NG��i4]��]�ݿK��T����c� )E@��Dc�o��-�,ؕOIH" �~�;���� �7��v����h�{H?|�������6	�6�6cR$���*6D­H�ѐnŒnoBf+�2���'�&�s:Უ�%/v�}k��?�d�n�AD�O�n��̻	W:,���kY�>��k��Щʕ"�Nt�Mf���t�,�B�����0�_��k����%Xw=�o
��ί�:F�iHhTjIY�j�P�V��D�7�����}��i7��$	��A����Q}:�ɘ�Ǆ~)��dDkv�0a�?VĨ��"c
�;Q����֍��hːq��"q�:�f������m�]��(�븤�F���u��e|zx����Ӑ��;8��7�i~#Ɇ`��A��E���*Ro"���2]l�6�u��q��L�_`Σ��>��*n/,}���(Esp���w篾Ҧ�������)08�ײ������[o�b8�4^Z,�a��lP��	 ��\"�×�ĥM�hZm����,A۰mT�����4�`���E)�q�!Nr��F��0;�ٿ~}0p�8��?M�\\��X�DW��>����W�JN��*CQ��w���&k��u�`�B�L�{�����Z5���k��R��%�ũka�(�@p��A8^�%f���B�G�Q�����9��-i������>!7%j{AG�S1B�b���&��� ���|�<�]&+�7����}EF��GI�G�z�M�����V'dj�Xi�,�C�޵�˿��ތ�;߻��z	B9d:�Z!G�/��]-�\��&�xZ��F�a�H�_m2'81x��
���V�חJmp��5lI��T��\>�R}��9�c���YF���K%o��}��f)sR�u,ϒ�I9��O������ �2�8w�ܺ���~�v�`N�x�̩��^��Ǜ��|��7U��c{���O��4(-M����t����!�Q��,ȓlɞ6��qTe2Sbo65d��xC��Z�˱]K�+x��P�m�"�zF�����B+��[��k��
W�SBc��*�"�9M(M��X,#F�n *%5J� �Z :�}��7���B�UȲ�*X2%β]��b�� h���<����]3�@{˦��G��<U�&�h���p
�9c�{ڔ_����2�l6�%\EQ��3�D�J��G!����S��b��D�/ �7��3~���o��ܒ~��Ö�W�f���Ty�1� �0��B�9��R�ϔn� �sY�r�mB����gՐ ;�㍖�ΎJ����Ű���p��3��oķ��l��שk�m�J����Gof��y�l�a��מ��톖 Ŀ������g����ҷQ��&�����-�귋��+Q�gD@j`������M��<U���S+������Fj[{���G�5�o�%��ۿK�*C�$�)�Y��#V'F��A�Y ���F�%|����47)rq����j�E�\<�@V����Uh�ށ��V��Q��O��V�]��ɵ~��ܤ��3"t	��٠>׹.�qJL������|�}-����a^5��M꡵�����Ӣ��u���� /�t��'߆���Vd�zX�Aa���B����(v��=�tkuق���?�p�;���imWN�y�4(,\j�'���f�f����c�L�ɂ7�
^X�^�4�`�Avp��DF����헁���7�� ���1�>(\�ݹa�r=q���v ~3��w�&��R?K��8m\���V~c���z?��s��='
��M�_�6�;��R=��l���Oq�;�eͿߕҠ��	08��q	aR2��e�f���G�"Z�ӂ=���yfO�����%��)Ac������ʮ�������, ��9�r��I %ՠ&�O�3���Ј��'"�hco��i\�4��G�z�ZN�ݯ'(���;^�1|+�`���%����b!��Fj�SL�;���*����	�����7SNI�G�]�����bLm�IԖ<��S�S��J�ޑ����ם���mf�2�eCGA5}����g�Tk��ױ���ۻL(��*����[t[-좬�R3�:HCE8�[k��"T��2r��u{��ć��)��q�3���B]�s[����x��-���M�o�p�HH�n�o�s��ki]���՝:�x����U�谥z���%�K1o|�u}@��t��/��-�,5�A�Gѧۖ4�C����
tW�N��9�јA fo��C����:rqkNe�g���o^(1���D�cˤ�W�;�.gJ�"c�q�G�h(\n�B�Vo�.Jپ��G�]kCv�B�Ă�H�'!pGJ��d�����z\�QpK��JНᤙ��Jug�:������c�XI�UӰ	�[���e,0��!<45 �Nq���1����,����6� �"�J��V�IX��Q���)�G�ֶzz|��*:�� �aɀ�:���p/�'�I��j�$���t6U"����p"�G=cl3��܏�>\�!�n��w�o&=#ylG�n���Xw�%@(�PX�K�d_S��7ίv2ʿ���%�Hq� ���s�zɿ���9o��_�#%z\%I>W��ZF(����j�=m�K9+bM�F���,�}WhƎ(W��% x�Y��0�)���$�z����_�-��_������c�w��l-�Id���zp�n�'��k `��x�@�ߘ0��(B~i��(�j��WȔkN�4��"`ɢ!B� $i��Ì;@�����!\�|g���b��U��.O��u��+���N�Ԡ���|�u
�y���M4>M�ʆ�d�v�~�G���`h��H��p<�t?�	J�N,Bz=6��W��TqH�`~|��@�FWa�w�OS�D�	��4�4f0i�-+�f�\���RӲ])Q+�k�`�+	��>7��Z��X}�i1���˧�DbS�ʛ���_��W�(N�S�߱���%-�Q�d�ŪW�:�Zhg	������7֟��@�
�Yp~�DЕjP�׬XZ��>�z�f�zW��E`��Ί���y�����::t���p0Ư=DpH���%:��}�s���9Avh���L�a+��ٮ6n7WC� 3%��~E.�t2��\��2�� ׺G�ّA��4�����.�c�g������n!���]3N-�<W�~~&(����p��2(�0�գ~;خ5Y*�j7�ok0�6�����$�XJ� 2�y�Ibj�n�H�r�N	aO!���QV���=�Hr�t^�Qu�:�M���ӧ$�HZ��{N�]n�x	��"^xC�|��+��O�z]\}�	����?��OS`d�x:?�����d7Ͳ�,��]97E��n���C��C��:wcF9�u�hi��z؋*YK:hi1f%��ز�-��R��h*{iW"A{n��豚����xo���sRSק���5���rI��H�
�ƕ�[�zu]�W�c�\�J�/B��%�q��[�B�̗��z�X,,͛�*����ii�8����Ģ^��j�q��B.�`�1��!�۴%RT��Ê��2 ��~��KC�#��\��I<����Y���E?y��[	uX�T�.�?�3�Q����Ǆ����q9I%��5�f^�όS���M��DQ�]_T�iS��P�̷��j���WsM�5
��4�u��8󇘽�]����*iC�.��=��k.ب���Iy���:�ߠ��ݡQ�y���c���%
O5b�\�׀��/�jۍ�%�y�ߩ�a��i���S�]���Q�<@b�LC���x��I9��|�:�a~ʰ��;u�s����R`]^���PSJ�x@�������m��s�O$
+8��A��4�`��@���ʙ��ظK�s�5�Rn$�n����h~�kdУ����{��~�!3%�2!�o&��FV_ns Z������!���c����'M���� �Oh�~n,�a;_g�Z��r��Gp��oA��%#��� �~��Z����&K�;��֮쵑 S��]�y�uc��i�ӈ|�;m����j*T�z�U�2���<-H����im	1�:�g�"1Yr)Ӏ��1�-2�_)� �-E�U!O7zY.^w�/)K<����Y�]ٌ.M�F.� v��u�ѓ�[7�]�3��kɓ��u�+
c���/kq6��
����Z��;-%@�.��	Q�ֹ۠W_�!Zd�l?F;i�ƹy�U���Nb���2�_+7��}g�fp�����+p���){�f��:�Z���eX�]��|!7�(�����+�+lC�&5�y�Y0|G�X)v���v �]N��៱�(����~ƃ�Qf�A���2��)A��,��Ja��^��7i��	�)-�?9`v��'�7띾���RŊ���c�����Ԑ��}@������pj�����{x1�Y0�D1�y��):ç��d��q_Dfh�d+�^Yh�/g��A�u!2�r�M��y�V#���>�0��m����ѽ����-&�u���*��x��I�jB(Xܚ����n;dQp��sH�&����#(U��v\�4	���m���1~0��v��hw��XhN��ş��"/�_r��u/�Ē�3��b��EgM�a��dM�2,���i��X�G^B���ޝ0!Ԏ�Gz~�z�'�M�Q�D�}2�J�#FUf�80��?�xa$�~�~V).@ ��dJ����<ٶ�L�������h�{]������s��R7��쭃��pU>�ĭ�>b��1pT#^Z�EYZ9�O��y��>�{r��<s)A�q�%/M�X?B��!��3>�&�Ls���h�?�H�Cؽ���%��e_��-��!����A�7� 3�-�]Hoo���BkQ�1���S_=�(�5���g��K�2�K��ՂQ�x\��.f>��+m����wG,�/���Ŕ7_V��31�3�Ũ�*��W�5l�{�N����b����i���H%���j�e%>zز+|�f"��w��r)T��p��'2%h�74(f�_��n����J�ѕٞ<{��"��I�f���E.��fp���g������t�^J����6�a+{t|�8h_[��S.}�����7EKV�p��絯N!,Ӻ�wñ�ݕ�U�˪��3�����}��O�^��@�*L?�~�j7�����(�:���%�Y�L|vf�F.����Q�eƪ?�=+����TP�`S�\=�P���J|'��mN� ��[A.A�X�(����;��[<X������x�\���*Au��"� 4�~�16	yE�#'��:�7#�O�C��W?x����<+��f;�����S�jif�/�
��S�z	׸8ÿ�֏d�c"hɞ�ڢ��+
.��.~��NR7�z���Z�}8%bɸ����u�s��(��Ά����ej��t��/ ��ҫ��2^�(�b��^�q-�tc�P�!:O��r�@�zG��ؙ��3�~䃒zp��:&)@�[��:�LS����{����TȇEe,�Ą�w��)}������/��͟~���������}�:S��J}���$*��F�J��?d�T�]�-LKq���S�]
�P�ݡ8���-�Z�]����Z܃��~���ެ�E��9{�����<	���`� u]v5Jh���m���"Y�Y�ra��(:��d�$Ƚ	�5�7�D��M/6�x���2@���zcj���K����G)�/Ǎ�*y��#.rȲ~��S�;ώ�9��ʼ���K��@1.sD���3-(��o��`c�DА{�?d��ۯ��	"��6��-�"
;8��=Q}�^'$&�HV)���eF]d�>��������Zm�*��B��~��F�Y�9a{~��Z�������P y��8���(��MPg�D�NC>j�80�.�@cQ�^���'����4�Z,�
*�kѥ�օ���9>_�\������m*����j ��m�c��#Ǐ4w��?����N˴4q��o�\�E�Wll�jG?	7�w�"Y�w��Qَ�I�[�f\f�Ϟi�=��g�u㐈���{���f65�~�	;<�V���w��������d[&Z�ߐƔQU��4#�(-��C���4�$��j��B�Y�8���4�� s�����+o��~��W:?t�������i>�&�c�/����e?Wϴ��~=�ǝ��NbS�G����g,�~1�v���H�ڡ� �vMG`�[)����q�+��7�����Nk:��j0�5����e�G\��Z�h,ߒt��]�(F��"�y��q��V��L' �!��d�.�����3K��� 3� k�%ȣ����ꉛ<��Ȓ�⊝��>�IRO�r�<g#c�-?��P4���Y���M�9������]��l\�Ÿ,��V�x�zHL�E^�~+����B,b#䌃&�1��Y�b�E�w��y������rLxU�%k�O��*�뒄�'�MfJ��h��Or|����Y��m	^��Y����Lu8��)q3}\ߦ[V���Þ�<����a�W�5�f�sVZ�$��ݹ�CZ��w(���W1������x� ��7AT�rlT����0�q��D�P"|u�~
P�ʻ@�6�q��o��J�H��p���k�C�v���5 ���s⢤@��)\��u-���O��H�[��SϠ�Zr�!u���xH��AV	^G����!j�ԃ(!C��l����w���:��o�y s�u}���\Hһ� Qi����sѵ��y�3���)^�g�o�/�B��4�W]�����$@N[�DsW�"�
CZ��r� $)��L�<R܊���~fƴ��AK��������:��[�}��`~�4����/s��-�����40y���W������2|���Uꬌ�G�:H]$G9�Y	���W(6����59�������G����j r��a�9&�_��W�-p���-	 ���X��[����7�/QZ�����%}F�����UW���Ţ�@uڤ��v�I�^q����V-�Br����F^`l8?����(e^4��d꙼���[�h�ɡ\�����y��]"|W+����c]�8�O[J��K_�梿��߬�?�BS����mty�AR���!�d���p*���0��-I�o��uJ!�0g��n�?-
Oz 9V}zy�CD`'��ܹ�@D/�����&�u������Q�]
Z�8��#%���ܬC�VI
$n�`U�X6�M���Qx��R�ʗL�d�̻��+=�񰳤?5��K=%����IR�Q
� *W�U�>%Ѣ!��%w�)�-З2O����]00ϕ�����P8��F?�EDEX��\�>S�+���wq�^���{�pё���٠��'�S���IĞJ��ZȜ_ix������b`���Jv>:R����P�axUJ��Gc��H�4�hiE/W�������C�[�25=A9G�^BF��/~GC���c��l[����r�|`H|y�c��h���T�ʹK�:8cM�;���5)��q%�9���3b��y��y����O�2�<�6�������=�{i���f�Thm!�9ou#�Kv�E;XQ�K�aEw�nS�K��Bv7��[��6o��.{	]L���<�|Ѳ�[��)D����뷣�	��Mn���n%���*���~%gQ��},'rƶ4S.���Y�͞�[񳙗hHV+Dh�ЫΡ���x'��(��.�'��Or��a@�[�NRiI�aJ��tȂʓ����;A�<��^+�1��A�[� ���H��#D�|��%�/Cl���.�� 
�n�5���{+!�����&mA�~����
��M���a��A�o-<۹J-�
�YҖ�� ��zg%�TAp�����s'x�R<h�5l��N�3H�L���Td�R�4���˛�J��o���`��V�;E�;^�b�������ؑ���-�/"�ɱ<[��v����I�8� 1�[�&a���xS���M�ŉ��OG��TiE?!1���x���0���E�j���nR�RC35J��� �Ț�-d��;�>z���~S��c�}r�iu>a?����vo�&j��~��AÖ<W��s�_4�S��6�q���n�L��H�^V�jq�#?ycW���MƵ6T"�:,N<�^~]�e���z�J�����A[ ��لqozt�W{�_@\ ��i�^Юn��N���dwoA�����8K����&d5�Jz�oLk��F�HS�zr4����4�m��4)��Z�}r��'ѱ����_'T�^�YO�ep6��r��{��Q����|�H�NE�P��q,5]|�娂��I��8<��x�X��Q�%c=���� ���h�le=�n�S���iEp�y��p�?G�yZ���[63�vy��M;�`�z��V�d�S$Ym^�W�.����AZb�;�h�k��Ԡ��M��O���L�n	��#\ӭg�t��$�����97��Pxę"�o��v�+?� Ь*1���tYZ^���
�]�����;u�Ǯ��`aAЇ��kz��.�+2���ӄ��޻
�G�9͠��8���7��|�F���QO�0�t=��ס4��.���x����]W
�%1<��F���=��ϋ�y���5�7������+ZS=���h�X�F�<<�%��f���[w-������K�Q(���e�NK���h�u�O��G�Ztg�-R�,R�Ń���ɴ�ʜ��Jw���bsީ*цN0��/K�kN}�
��l>�Sgm�т.u�`��5�W�BM7���Փ�|n�,YZ�&��8:r�qpbIX��V��F���6��O�z;+}"��ž���	ͅ���LћV��@wu:�$�4���[��}�f�D�w��ꆖ���zF'v=7� ��e^��)A�uX�v]��Y9�ڼ�� -�t������sK竬m�aq5놪V� 6� �2b��RaI:��_o_�jW.��1�A���U�Q8�*�P��Gw���[�����w��<����)ƉWJ0k�ׯ���{IB�g� ��hgQDY�13�A����uʛ�X�e�O���W�����8�F��c(���h/g5��e����3e�H@�Tcҧ���ע�����`�JV"V��E���9���>X�Y�4S}�A�0�_h���1�)��t�[:�o�K�)�bp��&2�g|n\�VW��b���B'�KX[{�Y?t��`��zǵm���|<��Ӓ5�r/#��6Я�e�!xÕ���x�	cFef�?_�y�u��?��O�l�#�-e��� s�Џ�v��=ז�Q����T���]���H]�,�Ǯ~?���>d��
J��\�o~��hp'L
W�
��[ ��v�ť�"S��\ -�9��� �N�^ςRn��3Y��`�02�`ba���,�1��V�����к�7m%ɹ�Ի�w߱��xH�����S����"_!�)�z%�5�#���Y��l�=�3�nz�jL� D�}\X�ˌ{Y�D�+����h��8Fy��������'��լ�g4Xs�������c2�����b����z�V��@�T�?�LW�´���v/y<���G�y�=\����\�,VC���J*\���[r碫�O��"���^B��t��D"��9Ok���ɟ%V�{�*?|}�P��;���;v'���
��T��_p0GvI�z�8N]d4����뎶�J=��66j<���:.�]�]�5�8#F"M.>� *�,L�7�;FԸ��=�&$���&a�9:�;��h&��%]��B����$$����jv\��F�J'��"Ύ�����%��k�uo�)���c�g9��p׀�S�z8e�Q4l�z��>�|���pl���B�� g��i�K�Z�%�у���y�zj0����;��͇�F��u|� -�΢m�c�ݬc�Aү��5-!������Y��lӚ}��{�aE�BC��ۯ�`Z�g�ou�+�=g9v��<V�l�Eg\�ܟ������g�q��X%=P.���_����o�`�+��Ɩ�%�ሥ��F6������V[��l��nI.T��2R��U�^�eObZ���N�|�5��e���i�m��W�g�W0�*�¥x���֎o�����NY���ك/�`@>c�uc��-x|Z�F{TX��VeS�.p.���R��}0��H�L�	���n ǌ�x`�ap����%�=x]�ٕ L�x:}�+a��4m5ˢ�ÓV�=��P���
�bS�]
X�DnU�0���9�r�L����Fol<�d�[<J!��}�I��0�����g��i�{}����ϵ� �4s ��~#x�|B��v�}�����8��#�k��	�%�Fy�j�-R��T��&�KZ�t��0�����P"��kTi0ź�Ǉ8��R1�� @$�[�n8����_�C��A5g��9d�X�z�E�P�!!�{3&&p;G���.q��̑��,��q���r��R�8{b��!DȍH�i���n���#�D��L#������k)�ȵ�����#Yt�6߈�<tH4�K�ƥY��cv����vy27���\�B�&G�N$���i�/-���u��{��U�~]���U�YYl[�t��Z��|n��2u��n.�p=�6u�tR��b�ݐ��~9���B�XB���l˕
��c�4�8~;gT�S�ծ��V﷐����7�녵��F?�Bc�2=N�s��&kv6(�Nɴ���>q}����Jf�:~R�D��IX*�����/��j������f"�J8p2�\q�l��)��D��;HÌ��@��9�f�0�;`֨��o�ʁ�~"c]|��\[9��U�B��v�GǪw��?
���3�or�!L}��X"᷺�
��ȑ�ᑽ�x\��N.����fU�(;�u�M�5��ɱ"O� ��� �nHW�5d		�M�)ROC��H�k=�N]l� *���!�f�+��P>Z����RyGj۳ż��GL)'���=�{т?�ڜf�{霛y#۟�Ei�m�Y��-x���	��K���l���I;���F�;6�����������Sw[���E�X+��I_�{
״����e�:
_gAa�ʴ����^�ŅC
��;�7������� �?@�r!�]?}Ü���Z��{�sӖYJ$����R����l%���6�T�o��������#��n2���C��X�U���w�A�@�k`ےі�3�����8�:[�~��5#���j1�@�y2����f��<:���:!���K��=�L��t�$��_�;���S��\�w
��mh�h'���k@K�
y猲k{��-R�0�L#���
�RT��إ����Zx1���W���0�s��{��`h��G�V���� �����K#F����}�d"���Ƿ��+�#5�jp�FO��ij�D?#�I�TZjDmӏ雛љ7.OsR�2��36ZN;���������4|���Ѓ�T	e��`a�OX%�%{!��H���ݘ�VP 4�C4*b
pvv��!�6��HJ�k�ކ۷�a������.n��<�LMp b"���xI�4jn5|	g�)����W;û�� ��nf���Z�JZ=��� ��Ot��C	#�Y +� ˨:WA�\ �)1��ZЊL�;�[P��/"���,ū묽��Yo�F2�?��6���ـlސ��t��M�:�'���y�'Q����z�X�]׶���� ��*�����S�KN� 7�'u�{H�֪<��*sXf!mw�M��{�������[]o���ĩ�d�5o#�!��4W7,�s=~c����a��$�2[�]�~�Gn$Y�wi[o��T<�ʵ2'��h��ZW����\���.�XW��+RG�Sʾj��Y��'`����e
MS	���Q�'�i��S�Ê�X�L#�yg��(n,O�V��(X�X��F�M����JRd[�E�i�V�i<�>�8�Cz^g���ml��ث�jm�Omtp���
=�=��h��C�m�鐔�C?�]`�> $e� ��*��x��Ar�W�j*�."=�k��Gg�#U��
a��Rn������YH��M��2�m�|����E�Ғ�7�V�ңL�@�}���O� ��q+�ΣUݯ�L¦��{[�}��U�n���}�Z�s�l�t�x�yb"{.쬵�Sʋ�]��I���0
��#�����̡�q�<!F5��8����AH�֞�ۤ,ިiX��Qy�v�m6��̀:#�l��L����$��q�9��
�ء��EZQx�<c�L�g��=D����|�l�3�R��H&,�vP��U�#ױxU��݅�9�%� �f5P��p�B�\b�>�@�cɩ�X;<��w*b�����,��P�_�D�hU^4�I�y��F۱ǣ�='�%��Z�m��K������ÝЊ�C�ԟK�Y�<����艴 ��Ⱦs��D�W�d	�#����Ǿ
ܫ)Xs=�8����J��9*8��M�D��DB�*Q��f���?�˜A�eg~�4~�Rӯ� ��b��������]����o�g ���P����L�kX)�Bs��ҖM�@�o�=�h*�x��Bce�ύ�j�-ݿ���e��LU���ڢ;��������v@�cLܜ��v�S=�������f3����:m�{ߨ^ƣ�0\3�dZ��<\t�v���p/�"��P&ɘHH�s$Ij��5��9Ue(C��kM ��paVA�g�)�����w�و�+R>Mfl���NHO����v	I�n�J���+z9������~�����3�%��,�O֚��ñ���g��L�>��]5;�`җoJ����h��ҩ�Vk��D�L�P7�{ϋ�i�n���t�P��ί��?�+�������h߳'G�V)}���?���'-JW���yDR�7�ɦU��˰dbd�����#�8?�-�}.3�y3�m��d�s!�~�6!�{ϼ<*���H�r폆{���P�~��3����"����H��yՎ=}Լ� O���YB�����ϸ�&�g�(\�����6?O&�apMM�*|�1_.>(h4~��0@2r��l��h� ���ǹ��^M��`�a�ڜUv����{]H��(ה"�:w̲b��~�уmD��&�]�/���_�c��{?����:p�嫻`��~�t��SCv�"Ay��n�CA�q	c��K�ʍ�w�������B-�sI�qij��!�AZY��ݼj��܍<���XL�}4�i��G�\�F*ٚ�r��)�Еv�HW��t�(Yiw7�]����V�l^ʼ�kh����sN.
��d�u;��:����a�_M��mH���w��I)�����Yx�#��!��x!��������Oc֣{���E<��F/��^f��т��nU<iKyZF�w,�.ey_D��<�<u�0��o���b���s��Q�;���j^D�v��/�78)`�� ��h�ŏ�܍5��}4mq�TFg����1lfI52��]���J<�]O�h�X�B=�5ʪEx���<c��Y��;�6O&<����-��d��P���[c��:Yͽ�b$�z ��'�&��z�
q�����֭/	�78x�p��5*H8;4yX!���H�|X�}�cg��&g=
T7�1;�)>ݰT�\�I1��hZ Hh:ހ��a�m�l�8K#�p�x��:���C�Uy�J�� ��`���O�ΣfF�E7��NᛦW�
�~v7Q��G�LM��B��}{���U���2z�u� ?`��Og���gp��M��ώ��Eg*u0����a��(���\�u�	���	x#v�;g.:&�����a�03"���BX�����S$�F��k������-�cF�N�C��5Doy=?}������RRi��Y�Z�u� 	B��� םa@�Ml�n�LxJ�1m9�^TQp<ޢ+��jcm���`1A=��?�y�VQ��|�3��|^`��}�Td���:]&0���W�
�h C��ib�9F��X�7�¿�_(�F�=۰�[R��L;�ڼ�nC�wo�#��#��ݴ6��f���QN��M��zr��V�:��)��!�ÍD-������$�6�/�$�K<�l���:��[,���nz�~��i��Er�R�b�z��I�sFٮ�54��2���8�#�[��K	��M��%��=�b|�z�-�J�1Q��F��=U[v�8��9�zY�����t��V`/�^�W��7��ӏ&����k7i��>�T�?�I3k�^�p*���+(�$=g��9Y���c=��~�[z�U��x�d�I2��B�~��y��匓M�GFA`d.��t��:�
�s��k���v��gA�Iw��M����z��w�ܴ������'>W���5�kA�NĲ�{؈�v��c����]Gm�BE���.	�B��,Q}��ܽT>*r�BǨ!��7��u��{���'s�A<Gn�״�R��D���_L�G��y�;	eD��)��uB+1
����CcR����O�PK�7L�k��Db��� ���  H �	��ms�i+B�Sܺ�G4�Z��^Kh��D{����G�Ʋ�ݙ�ŭ3:���Y�'��Ì�`zA �>rsR,�[��������U�C�͡��i���M⟓�Ք4��X�f┻��?l�R`4�C�l12��"4�g�� �H�Yz|��k��zۮV���U�B�/�-��jPa�Ң��:�4�@��?�3C1�}�ԛlnT�L���$�|�c�ѱ��Ħ��(��
ۭVa�ed>K�O�}|���]N.n�π���^�u��m'_�@æv$�~6K�W�|؄�k���=zm�0��e�5�I)z��>]�B<u�5>g%��k.O׫��<��h\�Vn[$�\��ӣ3zO��O9�\H^n<0�����
Z�	Z�d�����o��-�py���7'q����'�O$K�RS�對�Z�0zP����Ąx͗�����5v����t���f}9F��p�t�
�)d�s���t��tqW:�g��pl����B����e|LMH��N9�1���Xd�B�l���x�Y��1G\�� �꿚��R��&���G\~}���P�\�3�@%���l�����p0�t���hZǗ�����G8b��C<�0>0�'�k��Y��'�CU�Qa��O>��|����o���M=l:^���g|M�!*��6�9��OI�%������
�?cqȐ(������o���d]o<�h��V���6=�X�1�>6^��&�{������i�*	��T�`]������������}̞���eR-�@�Y&C�{v�+�_�\#��P�Xji��m��W�V+s�6r^sW.:�kN�<��z6h�o��D�}�X�W�,�ƥfz�]�;�t)��rI�!��DI�}y�m���H(�W�{85���M�kw����=[�������w�t�dI�517��*T�!��&E��O
�Oi�d�d��������D1_ƙ���w�~"�@�y<_�w�	lw��C�yko��ޑ����o3��>��G�G=�Q�q������i�V-|�Y��Y�(ՠ�QE�8�L��f��j��zy�5������'|�)����Mv�~�C�x˒#6Z���A(�ۿ���nYs:Ʒ?�<��=�������?�::�@��Q����D�r(ֆ3b	�H�m����-i��yտ��z��ҳ�[C�f˚�3h�I� ���)��@b\P�1&�$�V��{�v���S��g/·���'��@�C/����������n&�Z�Ów.=��>g��@�R��E]��n�(#N�=' �𦇪-�3�U���ߗ��E��@w|���2���y
��|�qwF�hݨN�����OR۹L��o?J3�h���r����}�j�z��QW�}bF20������/��jI}m;�s ���z��8�����񷕞r�|�#3�0�X���@A��`I�kQL�-�����q��FPqZ~"JUGm��R���x��G��������T�=U��o�E�~�]{%�c0�C2K�7�C��=���;r����[��p��_Р�F�ƒ�o���6�-�N߼������N	�%����5���bBˤ-��.�m��_�RM��1����r[ۆ-���RJ�U�*f;�_,��7ͼr��� �i�nON��t;�Ϙ��f+��3���|�_�2����D��D��
K�� Ōg�Mѩ/�ZOs��|+����cy[H��|�����'+g�:{��!�{���w��̧�O�ZV�8%o�q�B8� �D?����l�(�K"œ���(d� �s��4zT��v�b��CPm��9.�:��ox0��u�F�+��/��׺�<�e��g�'��7�OE�	�u�>�.��\Ԝ�<[�c�ƺ�P���0N����7�2�e6{�m�����@�� ���2��t�+�\S6���E�����g�C�9�\���!ӭ��.R�Q�Ё�{�\��C���$��y��b$���>�y
C% �̩��8�g/{��+޽��m�a¯j��{�O����2D�21�p��|R�j�C������V�\
�ot�98��e �]�puC��#s�`���
*�l����r>D��͆ �f��P�\��&�k��&��]zb(�wzXp����Aْ�,���$#�*Z��B����7]t�Ǹj>Z��[�sJa���-��9Gp���uWC9�+��R¯^
5NJ@��7o�A	�n`�e����֣y�N�<��=�����菓�8#GB;��]k��G��̟�9���87R����'��Cn�����Yʀ@�X~.b����q_�}Jk���QKs!gG���2�b���D�����	���.�h�xo��s���]�u�@k�h��t�B��ѩP���WX;Q��Ȓ)I���9#yɴ�mka�us�d�ϧ���`�2-�K�'��N����T<ש����H��M�:�?&�z��|��ם�4�S��d~���d��L�I�]���V�U�9?�Cuk�Qk���b�c�%��o6W�J�o�3yC�^��Wn��^�̘�Cfq����5�}&ts�S�}��Q��9~�|��Єt�@G�ĥ��5O���,~	CUs1[9�������C�/��?���GݍV�������GK*`5]�#=_˺M���kY�\����tN���	�m
�\�x,V(����~�}#j�t�q�@C[nM"NoG���֔&q(�q�ܹ
����"�_����۸%��wfvT�[���űl�/.>���Y �u�m�����뇃�G���p7�Oe����AG�z�w�s�j�w�5?�y:� �;E]���Q����S������E�W������}]#G�ͦc%���rw�h�����a�3�S��E�[,%mݟ��,|�fE�k�h	۵;	�z���S/�W���1���s���Q)�|,5y� �E������я<[j�p˯��oOܶ���q���EDAX7N�ن�]�tuR�qi%\R8�np{W�b�Z�"�oYA�D��,J���+��;�)�F>+�&��_��s�H�w��.�N�A�}��mF���������[�UX��D���w\g�q����L���ܜ���d␳�Z��Ā	c�qϟ���o�U}������x9w���dl�h�U��z096����/+b��������4�~�)�T9:�eOSe�Pz��v:��m*@`�����(���� /*�7�I�[)��D��C"��l���j�^�����S뭐V��3���<X�xO�I�I ���k�E�֡S{���6��;�*8�?PG�>>-°��1O8�s�Ō�lG�w�XJ�.���$�I����m`US�E��M��i�@u�o]j̰>-�'����&mMu�?�VF*�գ���黺�o�s��Z����,G��2k��B�t�t����V���؝:y;���:�nd��P	%��Q������V��~;&� ���FI�����!�` �Be�[Ԕ�h�U��q��6PeF��!L���A��S7gf�H��x���?�j܈���]����_�/#wWz�t=�5]82��>n��?���L7L�ֱT�(O�]1�
/�ᦳ	��x��Y�!yV�Y/
p1�[fs����>}���s\���g���	���p/�_���*��F�AI��D��d5DְJR����:�8�Mw���/����*���e8��4��]:�1T�(�ʿ ��1�Qȡgp+F[�"��,��b� �+(�8����#ݶ�_-�e�'�j��qRE2|k��?��F���<*�j�M7�+�����z/�����NO=
1�?Y��qf�H�2��i�lRca?')�t76�\�ls���Oυ��Ѯ��4���͏)T�..z�H����W��".k����|�RSdr+ǘ���sQ�$G�B}Xtr8[#+���!Q1վc�bbk��ʫ���ӅsNg��������.�2���w�*�K�(�*�W���_��d�RF��by̵S���VX�Ge~�<|�]�xe��E2�C{�'s2�#��@���S���ja���ԑÉ��J;�?���w��g'χ�Y�ֲ���g�c�f�0Q�3�������E�V���
,q	�% ��H\;MK�:����N�|�n��D۱��;̡A[\pbU��c�]	��z����R���ޓײ�"&��K�=��g���I�4.F���$D'�</m8�k�t�i��9?��p���P6��6���%����D���f����z��֌�Q��]"Έ�ݵ/���&[���ߚF�nG5���sd�ь��z`���՜0m�E�֍?ht(Tj|�b�6�d�y������2���G݊����d��L2���?1:�#�S�k�df��m2ۛ,�#C��>�f���[i�fO�m���@�>����>���B�{�b����U}߅�E>@[.�B�Ib3��:q��'��a�fb~xjV�Z��\�T<�ΐ��a��Zl?�2O�����'�-��r��{2���>T��>|�?�¹�q6}���|. Q��P.Hn&��!�輵��f/ަ&�2P�����k��ri�ގW�D���0s+sbSr�ϔLG�O�J�8A�Q2K ~gɡr�Vۼ�	��t)�����A�j$~��#w E���{�aX;�QZ�Aڀj"��?I����Q
�Ԍ�^�hi�;��Q?M���ͪ�^iڎ�6꾝�ѤΪ4r���ic�HY�:����������x&��\�ˠ��{��z.'d��묛�f��lZ6rQ���^:�(0�O�H�	Ӻ񷽦A�$�Ug�	���KWm��`vx���z�	7x�N�}besƘ���:��M�2T�0����k�7SB���e��]$�ƶG�Ƞ2M�dR7p۟�	�G�u|TK��e�ں]�L�2�
HNSp�ۈ���+���]�U���4�tm\�DO�E�;{��@3�B<��U[7�G١�E��nTj�Tk:[g�v0Q10�jO��t΁ɼ�V82�V��O�9rk��5/PN�6�/y�N�'�*1՚�������r��Q��ɡ��e���|�֫`y���uʵ�@�T,���<�@Nt�9,��K�"{1Lrhv����h6K�.�0�Mrdq�)�p$�M2G���f�>e�Rk��/D6���Mʱ�ǟ��:�%���B���I�4�)��gQ�Ć�B'���ozKН?
P�(�_�6��Sg�L�g)=�e<�����9u�ΰSK������<������v�z2N��"�>�~���`+��5�7�ă��">J��a�#KȈ�SN�`�����1G�8���"�ƫ�Ġ�x��J���ѷ���D:�K�n7��T?먛͏r9_���b w�w5��Y��Z	�*�/�=�7._�F}��Q��]#��@��+B�d���T�������Q(�oC������K�/�柕n��Ҟ�׹����r�eS�?E�{��VH�JY�>�k��O��#��O!�ՙ�Q'���W�������tc	-�� }nz�2�9Z�����Y�Q�k��\��A���c�n8֡*������ק\��mv�r����R�X����y�_۶��Xt3��e�5i��>[B�8g���=��$���:&�s�y������>Rf�q>n׺���v4鹜�qry�=?w��n3����C���_A��?���? Q�ɪ�6a�;��j`�Ϲ���i���~3m�wb %��:�L�L���
�}��A��1�����K�C`9�O��o�@7�����=
o7��a� _P)��\���r xܿ Q"�$��>n��Sm�I��U_rf�8���{^�IJ�G繜��9�C�t-�$҅��b����W��A)5����(�!Q��?T�2��^<���#�D���=Sʻ9��m
U������K��f�S�dO̎^x>bKA&��X��O��b��`D�@G�M����{�FɌ�L? ���7,�a��6Cg�A���(Ec֍w',k�՟�,;��Wl����[tW+ �O���3љ�w���U��F���)]�]�8<��&��/���@e7�I�����Z�Zk{��v6�E���q��|�h�h����ģ��U2 �MI�:XE'�+����_�)
��aASi1�;�K+K�sy��g0�L��6ѫ�����3;h,�j>��D��<E�{�UD����q�4&�� ��l�}<���#�&q/��>ř���P
�ܩ�'Ğ�I�+6@�W[b|�FR������Z�>h��q�g�񼯇�ߝ�����b��Ɯ�^uݔ�/����g�Yb�%E^���:�R�-J��
X���Rn}��`���oC��9��ʧlE���d��K�O}��6Q�r\�9�7�+��P��포�B�ܯ���N�X��	����l�G���P(����l�J�����!�l9���H���*�\>{k�q��H��}AK��"��r+��?�Ky1������W���+XAbDc�f�#���/��J�[�bu��y�G1i�J)���
�yε7�wВL��2�����֤H���Z\Pbm�ë��-�5n��+��U)��-��6'�㐸T�Z�M�]Ƙ�_+��n|�a_��V%���6W�x!�n�*B��J��g,l��Ѡ)�k}�wCM�Cdq���Й�1�w�\|���$E��џ>9��/:8r#7P�ę�{v��f+'.���1H<��'���2g#֖�R���.��J�M�yf��>�DaASN�k�`80����L4����c���b��R�(-o�p_� ~ۙ�hL�+�g��S`������E߾�c���Im�vL(�`��{���81�N4��0"�lJp]�.!���l[��T:mE��M0`�5�\�&��mY�f��������ʡ�7�L�ۣH�:9#6��?�X"p����r������DG�cR��Vdis$��]�&*B��N�ɨ����h��K��ą�i��K��ˏ�5K��!d�e��;���=�p	Y׬UZ:�����Z �Ҧx�ꭅ8c��:#V� ��eA�y����W�k��A�;���F��'@ܦW�Jؗ�u��O&B�:��t00R?KA��6�j������!x�u���d�	�Έ�%c��d���Ʉa�~�4gjB>$J^+�x�'?H����%�C��A�ߕ��Lx���W=�_Ģ������!��\�G)"���s�T�s�����2,���PH�5$��)��4e�?����R�.W�q�j૗�~�]q�?�;B�|_��῜�}h���R�3b�̺A�|�e�+�4@�Z-��bD]b�I�������p��E�a�%�v���QM_�@�]�7���1�B����QN/�����D�.EZ��X�X^�!8\,x���|��S�<� h�G��Y+j�����|��������3�� �
�Ɗco�(f�����`K������"����l�M	�2���)��'�=�&��Jԓ#bC^*&oO �>�W��X��\��U�k?��Ά��Lř�������K]&�9R-С�&!��_���	��#�L��s��b�����lCM���%��Fd%�v,���nT+*��4{	���W#N0�>�'ę�PQzK��|gTS�ҿ�r<�*�(��4!��t� ]��@h���j����J(J=�H�R��{'t�#�����?�k�_�e��v���<�L��<��|M֡�XV�����<A��6��|�D�U���i��iH��[����-�3H����ne\��/E\�e$����?��_��}|U��v6l�VH`�5�ז1�Ӧ�ݒ�j��6�QB|�� � L.�,S#��Q�v`w!�ZI��5��U4=�&���c��J�~$k���Ti���@K���~��O�{e��sR�-��(���-�$Gzk������^�iO�;�)��DR\i]��`f���,EB��'��g�=�Uh�����V��SQ9����y�X��@,�iD: �$p�����*0E�����j�(��h0oq�2Ъ�9�����qcrw6��9�L7�&�9\���]�������(# 侽Z׫FI��9�����7?�z֏fx�֝ �0��y �����)v-np�?�yGJ�i̒�=���`���!1a7X�F�í��*���>v�'$Bs�� �����$F���-/z�THl+���ϭ�T�N�@��&�\b�-����_6G�D���=>���)�5u�_9�#>d���0A���(�/�^���j���y[�%pH��y�Y�GR� B�{�,?V��3�C��X׼�P�r c�q8ޝ������(kJ����i��VHI������hw�9�Mb�>��l�jN�Cg[�`���$��\�J�3[����D)�!�ͳ��u�����fq���1+q����8�EN$>��<�ڞ� �u��{L�_=�-G��G�F�J��iih ��7��w�
ĥ��6K���~��Y-���ě�3,1|�w��$��*qI��;�&[��j(��H�y�9S$i�S��� w7P�Ա2��&'�����}�ei�q���w�W��{Vlڃ��Hb�z��]<r�D��H����; z]�����v�>L�%:f�6�`�kޕd=1l3U�����F���9P��Ʌ��(>G�ˉ�_��+6�"*�d.S�{Z�c?��_!�,x�绶��=�hH�bJ�I��/b�����5brʯ_��R�_AN*��Ai9ֹ���x���V�ON�;������~
��l�_��=�{�׊�J/c̸�[���Q�@Y���v�(m�ܴ�RI&<|3u�2�;c?Ѝ�Ş<��~>lU����Á٣"^�Ie�9�
lC������P�#L���*�s���O�^�-}�D��H�D��S�fyhM��v#�͙��e[���h6�j�N@(�e?�?���3�;���wF1�40_\sV�joe���׉ ���}��9�{���Y�~��I^�2���/��|+�����j����ҙ��w^�1ryO���b�]Ӵb~{�|�yƺ��&�l͹����.�q����6�`<�A,����B7�$�4�1DV�H�S[�)��(}M����f_.sq���Щ�K�6���;*�]ju�'�������0&ѓ6�g��?��ҵ֍I��k���b���j��9H�0��?�}*
#�Easn&��E�'k�m��vJ�/��yu���R-L|��%JK��h�'�3L�j��:����'�P�ӧ)�p��i��ީ�%o}2�t�|>e���:h�8u�e�O��בݩ�W%~��_ݵ}gl�9�@���,V�wVP�ӌ��B���Qߟ�sA�	�3V
�}T؋L�}��H���V�5g��5i��Իb��\D�<!�ǌ�.����Q��n�k�>�_>�u+ɢ���&z�����׾4�Go�p�S��+`��j{v�FoEx�
J���a���1��ԊL���!hk���m��޼���g�e��Q����齻���%d��^�	zb��fb���_�G�s>p
�$����ck��ɬm��ú
WV��
�&G��"2O�T1~JOfW5M��ΊSc*@O��7����bؓl�12<Ŏ�0����!O%|�Q3���7ν]N~�4r�CԄ
�(���<�
��!ZI�7����E�s
�Д�ɮ/�5Cc����<DAN�:��U$���B^��	�����9ܚ�����[�1!]�A5˝�-�Ԫ���!���<)�j��2�K9�q][��ػ�+�K>s��ïK�C!G��.��db�@��#+A<֨�[������s8l�,7|��p�͛�:���񮢼��Rc;�Q g-VO���	g��ᚾl@�ȎSg�N���qP����`�-�U2(��Bxn���^�ZB���w=�I�t����8(��F�Galu�Y��\�҅ ��bP�E.��3���?.[Ⱦ��h�n��E(��6�{�U3��V���:F���U���L^���;�����>"�xD$�݈�Z�gD����n�l�p[:J����у�^���*E徕�//:s�;HK��&���ļ���yy������y�m�/��Χ�PC[Wb�猯u������H�#�g�T�y�E�Y�ce��<>W��:��5�Y�қ�"_	�����g����n����8�n�nK󕼛��*x��Ss۝ �~n!Bz�מ�6��-f[����[^�s�� eM��MǼ:��r=��@��F��s�~���j2廬�M�7��E�|&x]]'V^�����`v�>�B���I���V)�����2���I6f�l4=g��7*4a�� �>*~⺼�H�pIM6�-iFm3�����]0[��).pA�u_GAAM��P&©�T||�kH-4=�:NE��8�H
296����Z=~����^7-��u�~>����m�ys[�� ��|2���E��+O��kq㥵����b�N�V_�&�˷�r�˴S֬��ļ��ng�����WE=�\�rݼ���6�ƻX���=�|��#���K�Yd~S���{[fl��AȤi��;4��� ���Ҋ�.����Y��-�f!�e�z��������Dw��+�V�6!�>�|��xW�ڞ���B�aޜ�a=&fEҾ%�w��H�N\�
q)�s83��U���<ٵz&���:�*&C� ��I��T���wW��t8"$DY69|+M��w�辯���?7q���cZB� �ķ���F	���᧪������x�EQ]ѓMz��U)爛t�B�6N?A�ֽL�`C���w�_-��EP�3E��N�]M�H�q"D����HI{��3w�@m���jF�$�6�ZJ �B�yx��-�Vi]�O�<S�~�k��]�.�I�+���e�_v�����z��f�Q&��{(뉡p�+�s�X�����H��B����j�"5��|Zk��$�=����+=��?`4l�k��"����=3Qx4�ܘ;��Fn&]f�V���Q/D��z~գl�S]ct��ڠ~:�h�s�l�ב�Mzѵ��W<HSUiW���.��aH��O&�0U߸qRk�SM&�i-�yxńY6��˜O�5!�Y���<�(����E-��=�~��ˡ�j��a�5�����ƩU ����U�:C}vaf�Z����U�e����(�TWTjm�*���"
j]kڐ#B�Ć�V3k�^��U��wbv[�R���UҦ���b^!܄�xL)7=��<Q`!��9�9���g���&��ز���u����(l~�I��Oj:�*q�-C�x��[����d�ƅ/o�sh�
��m�C��^*���yB�b�ʑ��ؼ�`��B�\���?*��8�o�:�vU���gy�)����x"ڋ!Mc$���.��V����<�v2�mF	p�9�'�f����э,�vj
W�����5�6*�����ٻ^D�ϢۣD���&S�Pz�)vz�dy==�����2�a�5����M�:�������p���Xt6N�3G�0������c�>!�UI)z�X�~��YNs!���86�]����$UtK��3���*������6�\���+`�xU3�UQ��#=->FnU͒i�I��z�c&�҂�i=	�[�����i�ڿO�f]Ii=K1�[�D�A2b���S�]���"��
f��a�����Fs&��E�9�/�!��]&�����d�J�=����V�����>G������r1P�E�x�A��za�����(f���0*�F0^��c������l�sE�Rm�������Z�ΈL� 0�e���!�*�>�&�N�BG3#߉:���F�4�ÖP>a;�L~iɔ��u�lhk�UtWN]jdcFsT�̚e��`٧
�i��}�Hk'�'�v�)�0o��=���ꅽ� �; �5��9A%�-�3��C��!��OMY���)��՘�oÄ'M1d���j�>0�vǡ�FV����'JJ�7^�d�K��Y��Ĳ�d~Ď���t��w)����e{�l�=���w��,D�N]��V�A����Co&~2�����d�%��r%]�9�_A��RZd�yv�L�w�|Z�?��u��f�BP"(�Tm�6yS�s�,�t�!f�� �^���e.�5�ɰ�/B6MW�>#N�ڟϷ�Q��+�MNoǐ�<�p���;w)9�T��%�y�%�w�`j8c����Y�SȔI;�ku���ܪdh��'!�l�L{���F�:�<������4\��v��E,�;�݅�Cx�./�)��.�����iu�����i-6��j_�;n��g��_>re�oJX�K�27Z=�u����7m��ڊrǂ2[��:�p����id���@�D.)���o0��ZX��q� l�bTJxs5�FN�1D~;ʜ`��j_'!n��y����XH����2��qO�к;VD9��]{zr��z����T�:9����t��M�a�:����r&�I&����Q�����up�r�o̠;�x�茪r͢}���3t& �縶��Eܕ .RW�\j7#no�\a��v��E�v�yr,�˒.8��*_?ɬ��厏zsಭE�؛�ͳ���<\D�f"�<$~z��N���y��_��Ȅ��/'�
�X�ŝ��G���Ε�B7zu�����q���� ���AG=��`ŪƟN���Z}з&b�ѕ���[ZY�4� �i��Ui7��b��SB����\���O7��6�%JZܲ`�������ycD^X�90퓺%��3��@u{=4��*#3mְ>����Gh����)�Kq�f���ex��k@��r�5�2�~���"�eI���L�E	d�|#E�vee��&�����:aj�s��[q[����S^U���B�bEN�V4�v�a��\T]�3�L�߈/�jh4�H�Zv`�X�G����2�q�-��b���<����c�l��:.���L�h��N���K�x�!��2-�:P�)�$r�ʺ�)*q	�mu��XM@n0�2M��ݍK�)�\���f��y��{uP)�� +�{�d(�q�n�Y�BT�c�.�	��2<���lz�-P�}�Y�
,�P�p�j��q����	BH;�P�N_o+w��2��(�0`�d'�9�**���f�9�U�I0���@N9r��
�������7�l!6aT�9����Bp�ԟ�
@q�|�i�L�OL1Z����H��ۢ�r��3{���]��ʖƬ#��g&�DA�V+�"��{��1�	o�(_����T7����(��#���L�c����Π�O����:��hs�\+�jZS���u�����?9d/F��<�j��h���D��U�_kDܪ�v���L(E�o���5���֐�<����\�0��k_�ݔ~�o�df��|c*��&Ҵ/�t��'����+��9��:�'�eEy���.`���x;�F���0N�wI���1RW�c�W4,����	R����kgZ����D*ՙ��fɻ��c��GX:�^�͹���}BT:v���@Q��Z	��gdϣ�q�[�2����\��+�}���W�~�<j�*��N�$�@ԑo'y�!X�l�m��Ê�q�@2�5�"�����+\�E�9"�� _�#y�N�F&C��Gt}orѰ���D-�r���l��-���<����'=�P�eq���>�K\���(�S|A�7D����"$5h\�h�z>�N��?��S���ʂ��������^�$,K�Nȹ <��/Y�<˥�4r_tg��(&���I�0qd���"���i�
��g�{"�b�o���C.޷�~d��$��3����}`MG{ &�E�25����Ĉԭ��M l�����	Z�g��.ўrd�r�Ϩ�Ѻ�gg�ý#-�M����w<:�}��Q-�b\?���w�K���d��m�R��YJk(��e6��k����KxH܎^8{���3�[�i8��%×Ff꙲T"��x޺f��M���3@���$�����0h2]�G��+�#���a�v���I��Yқ���D�q��!S}'{x�ی��th�-*�ś�w����g��@�y��V��BL�e����.B ����V��"x��˜��] �+*'�a��M���*�����#���s�c�A���Ğ�~u���Y�ۼ�1��"��Q�ǂ*0�`�H6��%� ��𲎔�N�����?��ap���)��P�}��	����|-u�� ue�%��I1=j:8�~v���[�~d�T�*槣�c�EPO���X�L�n$�*4Z��o쳎o?
Q�T��|HA���ˍ�oϥ~�g�;��2q/�������\�_Ey�������P8�s�bɻ�ĝ�)�0&B(�E�z�ü+��-/?"#�E���[5a��%�}ZZ+ e"Doq�g���'Rm�U��*�����U�Gb$X	� �>�͔S;Y�`$��U祿��r <A�r2��u������#��̇9��W{���"�K`.Xfa[�U'ٜ��R��bh<��{���
R���*�* �L?>]��L:�Oy���Ot�^►1��b&(��*=G�6����2^~��s�VM������K�1�X�����|��0X��9�Ogz��@!ޜ�0IJ������M���u�}['h��ow&�_�hO�)��F�_�d��
r|k���O8ߪ����CF[�E�	�J���!��ʕ��Ǝ�/ɽ�������ukך�i���b,� ղ�pkB����?���x�tu�DЭW�PH��1'������S�R�$xxU(O|W�Ş��Db#i�����<���^,���Bo�"���HuA�2���#�i��F-YC�!���K}�.+A��P&¦�����)!'�ȡ>s�'9��ݥ�jNsO��QcC��5�eI�pO�◱�6���Q���`��	�rLaM���m�Ԁ��%��lw��Z��c)ϕ���y
L��h.7yz��Q*ɍ��S��Q��l�}�XIe��Y���ɩM ��i�e%�4�y�_���	r��LE��E��!j0���ɲ��)��S������`׆�Ǳ2ޥ������d�,��[��.�窘�J��7�߽���N#eRǢ��ɳ�8��>���	z�q0@}����j]��l�t>�)!_(VX	ݺv��V�4E[�N������3 �������$_�.��"j�����Jd6^��&�~�I���I8�H@$GT�&�bˆ�Id̲(6]����3m�[�,(,I4a������DT�k�?�\J���=��(�K%�:Y�H3�u2r}��h�׼
Q��u��m� �82"����%��L���%M�����Ċ8T��Ha}���[U�dX�>.�6+��'��tN�ʖO�ٰ�4��ƹ�NJsEa��/��~&��W�������L���zD�!�-i��1?�c7o�aR���:�SGg���pY��C+߰N��4���m����CZ'��N�I܏�_��4�i�C�"�a��Ä�$��Оqn���Yg�m��Z�̺�����'�{�V�+��f���{.M�7ʷ�G���135}^+��B�z��o��ڠ�Bo2g{�>jwb$��Q'�̐��p �7j��PX���[p��r�Aw�5e��M��W'���������b�1�n)^[F7��x ��:�����/iڰ������k�o����A-�\��Ǳ��؋�;�ͷ�pK��z/{wk�N!���V��Ҹ��u)i�x!m�������A_�F!s����?�?���_����G�/9S���ҭ'���8�������N���H1���?\��7�s?�$��_a�}T�����\b�l�255��7f��
`y^�N~��g#�m��r��|�;]mdĠ��myy�����NNN+�!��1��k+�h�����Pt��eT5���P�/���b���/��?�1m���������_�/���b���/���O���˿p��RCE[9�����PK   �?X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   �?XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   �?X�V��  �     jsons/user_defined.jsonŗ�n�8�_%��4xE�;m�� n�)����D�Rtiy��$���D�n�N�ȏ���?�c��E�ֺ���43:	f�]�Ya�8�sd[�6�������˅�wc�U�f�8�����l�mQ=ڎ��LU�*LSy���f�O�>̳He^�Y��� �$f���S���8QLlg�R��Zת��f���L����$�,Dqh��X��:Ԋb�$���֎K�� �5,�jњ�~(3�1i,����Y]��qU�u��3����x���0pإ�d����l�mSev:��]��κ��d�mA���݇�^uWTvH�h��nM.c�����ޞ����4��t{����������X慽ҵn�X2Ɔ^X2';'���܋��L6fF^̏���ⷡ|����m.h4�b/�:�b�t(�-���XV���/�:�;�K↎%�������cAa���dn�XOB���B���nꄢ�'v�tc'4����c �
a?�1�����îё�5���X��D�b�X�h�D�
}���O$-�n�DΊ<���:�Xk�P��:�F���MK�O>T�-�'��/D<���'�-/<���'խ.2��BO�[\d"yqO���M_�~��CV�b�َ���P`���4"��Q@I���D����K�B�C�]VE��&;X��ߨ�@m=x�}i:�!�w6Jvή�9�w�åY��gĝ��eu��g[���>޾���5�4m*U�V֘�k������*;�0�4�?��.���\X�4���>�ߕTw����5W�V`{��u�T�.L�ζ��E��jmL�6G�DB� �� A��H&(�%D�������4@4f��#�
��B�F��4L���?��sF9��Rb�!�tC�1����#���;�j�Z�ૢ�CN��7r�z��x����aϧ$����W�.OqZ�_ b���~o�����~E���`]d(�uoKY���5Fޯ�a�C-��)�(M��XA�bD`ɃN�n��PK
   �?Xu�ŋ  s#                  cirkitFile.jsonPK
   �?X����H   C   /             K  images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngPK
   �?X��) oj /             �<  images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngPK
   �?X$7h�!  �!  /             Jf images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   �?XP��/�  ǽ  /             �� images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   �?X�V��  �               �: jsons/user_defined.jsonPK      �  ?   