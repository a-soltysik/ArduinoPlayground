PK   �	DX�v{,�'  L�    cirkitFile.json�͒�ȑ�_EƱ�%���uS��t�Q�hL{�j���mv���TK[�4/�ϴ�`feA�������}P������#���/�C���a����߆��n���H�n�S{�i���ܭ>���������O��_����?>Ewھ��s֡6�����4U_����m��p�֑u���~m�f����o��̚�Rfm�Rf��l�����_�Cqhw���?��������a��Jv;^|;^x;��v>���ķ�n�O��B)����6��?�������CŖ��֗E]�Cai0�k�@�\[/����0�*�R�o�='�o��R��7`b�Є��0�7bb�Bތ�ŵ�5�[.�; ��+
�;0�;��U$j���ށ��"isE�D��j�����M�؄�E,>�m���ab����BކYy&6a��,�����Dl"R����H!��b�B���&"�<w�M����N��H!ϝb�B�;�&"`K�;�<w�MD
y�t���=&f@���<��~�{�ф� ��N�3gd���[��H!o�&���[��HA�Y��NWހ�1���/l ���	GxG��"���&��H!oL�&"��9���.6)�)\l¬�<��MD
�@���9=Xј�lD�N�ށ\\�MD
هi6 �y{ _���A��b�B��MD
y{ 6)��؄Y���@l"R�y�&"��_��X���y���!
�9��QJ��&�|�b���vº=�{����O��1��X�[�ۡt��3k�����J�̟N�&����z>�iNa���[�5a=�����.�o��+�����ά+��*��t�T\Y�����z��zJGX:�n��k�������?�X�a������CK*(��x�9�`m��#0O�����|���`��U���|�P �?�V�����)���+X>�d���	�De�Lf����j
����˗�>�Z:��>�>X>�����<X�`���K~���,��x���/C�OC`�c��ǂ����|�@�?����������V?X>��<�����G`>^N�X�`���!���,��x	'�`���#0/>On�,��x�,�`���#0/���?�|���`��g���������X>�/͆�/��K�7�l�2�o�.ܞ�]`�����G`�t�0ܤs�X�����q?X�8���������V?X>�q���<X�`���%"���,���B�`���#0_ZC�|��:p8���������@,��|\��?��,����
�`���#0���,_�|��7`������|\��?�|�����a����G`������H�}`������`����G`>�$�X�`�̗�������8�����v��]d ]e �~X�����������V?X>�qy7�����G`>.L�X�`���%���+���G`>.8��yݕJ�26ȳ �k�9乂eU����N�	}�h�{M=��ma9�i�ϥ[��N�V�\x��\��R��������/e$��O��]����K+I�}Z�w� }��/S�A���S�7���U���/��dWʥ�OkJ/�VS�辔D��O���Aty�^ދ.o��w��;��k�ս�������K���Ɇ��7��[���=���?�lQ�ޖ�O]��4�hK[��z���U�+=ЬӅW�o3�N�o2�N�o1�N�q�N�o�N�m�N�k�N��免4�qw���w�0�t��Ο���M�7���Y˕E��6��ކ�C��W����罟u��S?x�b3l��/뺨۶/��|g+�޵�RV����-76�MQ�{[tLAu�Z��_�z��«ϻ.�����Xߘm��v3İ��)l�]Qv������r�Y�����x���_o������I��V�b�Vw�7D(C�Mb�@���d�pb�FCT7���ˈ<�h4�?�}PD'C�ߴ$#*QD���v�ʈ*Q���E�l�� #jPD Cf���R$.k��6,o,q�,���b-5ԛM'd�%�K�0,}�,m���!,��,5��
�`)�d	��,��,!���q�%3Y�:��<nayeɌ�� &X��<��d�qpȒG�AL Kfq1�,�q��d�/ &�%3~m 1���q�%3~� 1���q�%.�c��q��(K\�
�P}:��ϖ c<���?�`ye�K���`y���8��8%���`L-R��l	���(Kc���Bϖ L�AqX��<����%`L�����q�%�� c��q��(K�^������S���pʾdLY	�`y<���(K�fԳ�����	����Q�x�)�	��,��,�*I,���<���k�`L�<^���s����.�[��!��
k�����rLlb�:]j��@ʚ��"�0V��.��[�U��TX�zZ�n�WV�����"6�NK�`<��"�k���uZ��WVRa�}�NK�`<��J*�f=-��
��+]`E��i��_��r0�`%V��ρ[�U��TXyN��0�Q\*��C�s�u|���4hI���h��VGy�В-�5���R�%Z�3��[�BK:�<�_Ƿ:*L��thy��ou��
-���Z�ꨱ���YZ^S��[E�BK�h!�tD�2Zҡ�5>:tt�
-���Z%���2Zҡ�5W:�U�"��ILG�Y]fut�
-���8���2Zҡ�|:���e*��C�ku|���ThI���V��VG��В-���.S�%Z^��[]�BK:��fWgb��.S�%Z^{��[]�BK:���ZǷ:�L��thy-��o�f+*MW��eNG�9]�BK:��6_Ƿ�ґ�6�-]��8AG�9]�BK:�\+A�ԹY�out�
-�|Љ[]�BK:�\�BǷ:�L��th���o��.S�%Z�%��[]�BK:�\EǷ:�L��th���J?����h�H�*-$SZI���Th�֎�ou���В-���.S�%Z�}��[]�BK:�\�IǷ:�L��th���out�
-��rM-�]�BK:�\L�tt�Z�Y�outY��e*��C˵�t|���ThI��k���]v�m�[�"JU>��|�負�˂�.S�%Z�e��[]�BK:�\�QǷ:�L��th����out�
-��r�Lߖ:�L��th�֧J���e*��C�5Ku�6U:�9K*��G��Gt���5��-�M�/�����`l׶�l9��B+3�iZ��&���L�Vfjx/�2�w�B+3խZ��G���XA:�_d�����K������u�L��mҺ��L���f0!<�{�R33eЗ��8ݕui��8�pv���(�����6�K�<G�t?�f��7ӭ˗��D����K�`�xn�ĥfN�8��ci����s����>t�-㟺:��4�hK[��z���U�۽�,+���B����B����B���oS���/S����R����R�������/&zo�j��`��v�&������~�)\h��\Y��o�,�m�0t}};�dY������~L�އ���m�˺.�틾!�ي�wmF�̱r�J[nl���-�l���)��\뢽���,YV0,7��e��;���1�*��v3��C�5ۮ(�M��M����K���~�u4�>�׏��8�>~y5�|{�{�����-���e@�N�
!2c<A�@���"�!3�U D Cf��@�@��؇����?!2c�B2d�~"�dȜ�����ڸ���K�(K�Ե�0�r7��7ʒ9u�1L��M���dN��&X'XGY2��_,�[XGY2��i�������q�%s�0���q�%s�2�a��q��(K��������Q���k
F����q�%�Cc���R`y���8�׋�1���q�%�Oc��q��(K\�����Q���
�	��=,��,q�nL7(����Q��.�	��=,��,q ,�{XGY�u�O?�<`ye��9Ø`y<��8����1�n�>o��x��q�%^�c��� ��(K�����%,��,��.,���<>gi�Z�d- ��iI�*���
�Y'� �V�~�`%V�N� �����J*�f��eA[�U��TX��R�kR��VRa�� �&�X �`%��GQ�kR��VRa5��*Я���j�I�U�_5XI�լ��+h�@�j��
+�	�:�K��thyn��o�T�����]�#�HGy�В-�5���R�%Z�3��[�BK:�<�_Ƿ:*L��thy��ou��
-���Z��1Zҡ�5%:��Qd*��C�kct|���ThI�����|X��e*��C�k�t|���ThI���\��V鋘�'1]fut���e*��C�k�t|���ThI������VG��В-�I��.S�%Z^[��[]�BK:��FTǷ:�L��thy���out�
-���]��I:�L��thy�out�
-���j���2Zҡ��:�U���4]QG�9]�tt�
-����|���2Zҡ�:���e*��C˵t|���ThI��k>��VG��В-׮��.S�%Z����[���ThI��k���VG��В-�D��.S�%Z���[]�BK:�\�FǷJ+ɔ����2��˼�.S�%Z���[]�BK:�\�HǷ:�L��th����out�
-��r-*���2Zҡ�Z*�:�L��th�6��out�
-��r�3���2Zҡ�Zm:���e*��C�5�t|���ThI��k���V�ʇR�]ttY��e*��C˵u|���ThI��k2��VG��В-ז��.S�%Z�����RG��В-����.S�%Z�Y��[]�BKy��[E�]�Zc�ؒ������~(,�vmȖs�0/�2S�v���j�����^he���B+3��Z��n���L=�Vf*H/�2S�yiԁ��s��.5��߹�U���D���K�`bxn�Хf0Q<��R3����]*���D��^�K�`�xn�ťf0Q<����V�s����>t�-㟺:��4�hK[��z���U�۽�,+��/T����S����S���oS���/S����R����R���oR^ԁ���{5yf0�{�W�g�f�Poz��.4uTd�,Z߷Q��6m����e���|NYVn?&��C_l���e]u��Eߐ�lE޻6#o�X�yG�-76�MQ��^�EG�TW�u�^K�m�,+���Ͳr��Xߘm��b�ڡ�mW�ݦ���tCen�%��[��z�������a�����H�n���0<�?�G+�z���������}��f��?��p<�����zr��{\�_�	'^�+�B>6������qk!��u���3!ɼ��B�֢�N��R^�=��3�,x��,�8A�����]��J�������Nzu�e/ʴ��o�$zq�z�RI������e#���{��I|y'���^����	�{0����/��0���[T^�CI�������߿����1�
-�1TR��M��TNH��@�[� DmADJqR��.�!L`}��Z�c��jB��v�@H%<��sT����A:9
�KQm�PI0ұ�tC!���C�ze��"����x����~�xl�������o�������Ӯ_}�"F��}-k��&N��bf�� ��0��	!�0��42(/��	T�C��ɠJ9T�ByT%��(keP��N=%�%f��(��0�ّ҄��ˈ���H�r�4�SʑfgKB,@z�4?[a~&@��Zؖ EӅ]� I��,}�)߁H�t!O�B,@���0�uM�N# S[@���0��UR@���L-�aNk��b�8L�!�aN�ˤb�<M�!�aN�ۤb�@N�ȧ�O�6�i����O ��m�~M @>u�|*��� ��BM� ��]��
E ۺ}[�nr��+���� 8 ������8�(�E �LJ� �Xnc�̔�G4@H'�R,� 1 5{@j���� @W�����cp ��d[�.��~ȶ�B����ɤ˦X���LJ� a��q�r�Qw�N&�X��r�� �Wn���8 �7 ����'p �o	H�r<%�ȶ%�o��X>Y5����w*&)�G`�d�z�҅3���Bw&uO����Mn_:S�k�I�S�=�;�|�3�d�	�=���|�ʉ볲ޱ*	��dg	��'|���Dg���ĝX>��>�Ɇ�����Ϭ��!p� ���%��/\~��vBw&�@o�G`>�N�|�ك��G`>�ĉ�|����Є<�C�����'Ϣ}��-`BB��_���LHhB����!Z��		M�S��>D�0!�	y�7ڇh�&$4�IVCb|�N�k�1.E���y�Kъ%%�<�R���!����8�Ǽ�*LHhB^���!Zŀ		M�K�>�|�}A��V1�b���&�=h�U��Є�	�C����R�}�V1`BB�"0��*LHhB^���!Z��		Mȋ��>D�0!�	y� zn	Z��		Mȋ�>D�0!�	y�&ڇh�&$4!/6E�>Q>S�SZ�8�N��r.Ƈ�
�x����. K=��--[���&L�L__-��q)Zŀ	y%8:,�*LHhB^Ŏ�!Zŀ		M�+��>�h&$4!W@��b���&�Rh�U��Є�1�k6��c\�5`B.1�K����ry��_���&��h�U��Є\��C�l��K��}��-`BBr9�ѲLHhB.e�a@�0!�	ӝ-����Ǹ�b��\B�h&$4!�;B�-[���&L���^�If�R��r�)tX�W�×�UL@���V1`BBr}/��*LHhB�M��!Zŀ		M�u��>D�0!�	�&؇%Zŀ		M�n�tu�K�J���&4����(M$�����	��txᦠIMǥ�
�Oj(.<?)-�x���E��K�80��c����O*�.<?���H��M
�.6q�J�5�Uo�i����-5��^j@���oK$�y�o�}}?��n_߶o����w'\�	��M�o%}}'ҥ�.�+�z\��[KHc<��j��4���/mi��7��� ���m�������E[ڪ(��֛Ά��^�d�/���ܟu��ԟu��̟u���"��+�D��W^���Y�_�~�ŏ8 �x���g@�׺y�Da����M�BSGA�ʢ�}UQo�І���kY ��+� ��k�������a�-|Y�Eݶ}�7�;[������rο�_�rcC��lɷEG�TW�u�RK���g�/���e�%�7�7f[E�n��v(�f�e�i:�)�P�k��u����[�������:�j��*�1\}�a�:�q�̪�;<܉���!�N�X7z\�0��7�{Gc�k,4Vw{�c�s�+������3,�a��gX>����p|Fl��2�b~�\�;w~9f�xQ^O�'�DVzS�Ĝ�xs�O�hx���c43重�|�w�a�|���P8�w�I6%�RBIg8�4)�y�$�/ y)��=���0��s��)n)�MGߡ�R�J�kf��xX4���p�\<��5�7�֢'�H#�#YBkQvNv�H�d�Ǹ���ݘ.�L	e�Ǹ���0�zƲ��g���9e��(1�	S�RD�-��[���+�^~j)��҅�Iӯl0ڤDV�pe��t�H�bI�%��O-�D_`�Is��͛L{#��ߏ����Y#��?�����cI9�����'���Mr�?��'���O
�?������2��z��J���ӟ�矚�'z���H�A/���!��J=B/��%�rߔ�8��8�wN/wN��˭Sz����mz�����{yt�>;�5N,�a����7���a�_�����dEy��v����!�˭���C�_���o�<��e�������p����ϟ�_����|<v,[ڟ���׻����'��߳;J~�O�H������/z�o���㶽⏏��/��]w?|��a��O��Я>#ft����Ӷ�������ސ����@Qb�;���?ֹ�o^��w����C]˴�&V��]��U����mL�Eݹ��*T�����Q�e8<���������>lN���@�V��.ZiO����l{w��Ϗ8�A��w�w|;�9�����s���s��;���s��s��94����Vϝ2}|_sg��3�)�k���м�Ǐ^kh����y��|9	��M�g�2�@�i��L�T�ZL�b�@�<���x�90����v��4�.������мp܏cN�_�㟏O�n�5���`b&m���Bз������?>�O|���o�v����'��]�W�yo�S3Q�m[��m�.uQ�\^l��Ի�k�ؔWv���n�>)�4�C�.�'��Ű�M�P�rs3�M�n�8[�G6뺶9�g玫3�|�o��;.ؼ��Ğ�;�����y�r�@n��,r˜w`i3/�3����������}<�������&'��7�3���u��_^~	���2��l@��������w��?46D�|���t_��Cw��6TE���"��uhM6��"+d}��H4���Wŝ7 ��y��&�ބ��&f�Q�RY>ȇ����5歽'��n�}h�����,�"k��_.���R�䢭���u�Mɟ�C���F��n��o����s
���r��;k/���z��7��A��^�Fux_cjw�=��[׷���o嶰]�æ���Z�j����&k�DF�818��t�����?��9���O�d�������5y���Ou<{��G���h�s�SQӮ���i��	�s?n6�G�"�=o6�;��|�ӿ������9���׼�n��O?w��w�������7=����w�{Z�1�I?�[�MB(c��u��1��Іb ����ԛ�f�Y���a�ן�3Y4؉��h��4��Ͱ�������G���&|0��9��?���o����O�ǯ_���0��^�����8������OC���!��������_�g|tc~�]|�?|Z}����?��O�����k{8~�{�c?�$�5���3�Fۇ��?��-��"�}��̋����y�{8~�����ӊGe��������=�_?������-֡<58����G�vzԏ�~Z���[����V���� 8���r�Ė���`����}���z��]��ˬ<9�]<ʾ�K�*�l<��a��هUy����<�C�_k|�N�ԋ<Ok���=�G�y�B�R�PuRYGY�ɘy�a�5�as��9�L�U�1�o�.�/:ks�3��r�3�����xj30��η����"毳Gm.���Q��2�x�76 ��<2 ��77���G� �K��C��Y�ޅ
|�h>���M����f:>�19�M�.y�ϲ��.T`��3�d��|�L���(�y�a�����q���{��|x0]@_L�\Ǻ�r0M��w��>�o3��ׁ?~�0�8m%��w�;T����t�VK�����������G:��4}��7l �o� � � �4 LV ��
֙���oZ�������z�<�J��h*��iq��y-���b��\�d䫋�t6�>��$X/��v;c�aX?�x��)b�Ǻ8�l^Ocr�Y����sXA沺9�'�\�W�f�j����Q3/�W���j������J��]�d��bT
! �
OX͇@����&��Zt [!R�v���f��5�`:�:����˽��>���z��ug��e6A�m�*��.t �����p�v6�&�]��,>��������e�/	���ϵQ��.C����`����J��Л.�����w�l��|�l�q����7��׾B,�g��7�;�vq ڬ�7=��������3`�w������5z�wS�uq�5y�orX9�)�>���yXq>����9�y��3��ҳ�F�
����1��͛��qv����[{���w���8�������O��w���x~~d�]��� PK   �	DXG�~��  � /   images/0739a1b1-a163-452a-a325-ab452d55b136.png�y8�m?�r�J�M!*IY��Ie�^Y&������[�d�cb�0��d�1̒,�ٲ�L������������|�|�4}��>�r}��|��mn$�_l��mۄ�o^�ܶM�i۶]&{w-�����A���{����� ��n�m�&�I����em4�6�l����
�*y�����x(����WŶm;����5��9t4Gb&��Ȳѹ�}��OܜΉSٱ������b��MT�}�L�1HƸD���?j��i͘�ǰf�	�A��{�ξ�[_����J�z���r���٢w��/5a��t�I��ե�EnhǶ-?����'m�ں-��Ǔ[�n�-��v<����xN��J�h���e3��2������7��=V��)u!";G?�� ��<�|K0�yY���I2,���^)�Ϭ���Ev�p�����������d���4���dK;!-�L�^�$Cx�䐦W��k��E���9謗	* P��ϕ�����S�����0C���~�?��$Ǖ���φ%mXJ����{���w/�y|
�T!��;��G����쳄�[�����⩧�U�6}3���6��{�[$��ab1�P��~z�3������Y�q(�V�f��¦�&	�� ��l.Z��s9�2SH�W�ơP6�[��SnT�QokF!s�Ǔ`��� 6rl�������fI�:�v�K�|l��%����)�m����}gw0�6=y�dk��?�/������<�w�}l��جJ���s�+����������6����Í�͍{3�����"R-33�	a\yoU+����̡-�߶~�S���v�ѯ�f��nY7�߼�K�pE߬�����f�J�\t���+"D�,�����AGf�H��X��i���&���oց���A{10�^���l����UL&0���ٵ?���E�)�Q�5��s�=[�,�8�v�Y����>\��>\+sS�N��88y��</�!-Ot�HS�/'9��q�ZwuR��
���ӝ�v�����xS>edf5�Ի`��Z��/�j�3�QM�/
�1Q �wH����G�h�p���"[�|���fi�h.��-
��f�:�[<?>gh8)�2d����q���j�GZl��Ϩ�4.{��F���Hq���5�1͸�m2�2~�l����]I���J�&k�-�x�T�/�O�z�5�k����8��JdX��a9�<��V��\�����R��9�����0�TƦ%r�hm�[o���b�Pԓ��YپQ5Y�� �>[Զ�f�UG~����bhA�A	���6��,-��:[��Y����p���m���k���A��p�ʂ�K��&�{sdJ;?=3�O�	}�Ij�>>wE�Ws20NJ]=X�uq�g�j����bN���|�G����Q�s˪�r���W��ӕ������7�[����v�ЂF�K^��FY�{��s��ʻ��R�:i��D{��x�����T�Dr��j�M�s3�����:u˙��[�.�[Im}�v8��0��d�Y�S�ܷ�BW�V�F��V�E��V�
���355;����҈�RW&/�+�'��]W�e����v�@$�Y��=�Vܲܽ��ٳ�6�tinb��[s!ޞ�C����<_��iG�Gn���_a+*�� ]>��-u��{\lrǹ��x�|�b�ߕ��?e��@�㕸�����[�`J�p-��i��m�'���n��:l�xm�pd�l�em,W0Q�:��"�A�fXDyP��pOTG^uPiN��c��+l����~ŭdyώ�ȂrZ�����?���A�Xc|O���/�Pc���>���tx/��g�N8^xai=���
\�ΟNXi��@�l��]Q�0��!a�+ץ���q�����`Vq,�o"�B8a�i���Itq�����1C�06�J��J���
�<-VTy�����kQ
�ɍ������p�F����Ϝ����r�}��O��u�~�Ar�u�����Wc~2�ƪ����@�m�����
&�H�;7��.2g�>)l!�(�|�v�z��[�TJ�й��#�J�:F���R���:oȼ�>33�w��vå"����P|�?{�&��#�H��+���#��<o��Jڐ(-�������&�Mt^��R��|٢����q`�g��c��j��02���)����F�;W������+�xR��:P��/�ސc�H���\k�Ý�/���d�����^� u �Ƚ���c��������-6yK�.�d�j��܉�x�������7�.{��"�'�>����K�۰o�g����m%���UY�> �/��
zo��X{_�v��Kû��q��Ŧ�ү2#G�_Z&�k3��x��r��2#zל���@�[��װ��^_�L�#/=lql�X4Xm������nq�p�7ME]�A��J60��e��ogU.Ė�FՄ�W_Ћ�[cT���l�hze< &��x����/{�"�Lv��
��= з$:��Ln�_�|_�!��ɬK{U���G��Jak�6����������R3Ć��S�ۿE$��|��ӝ1��E}��q[s<w�R��.�$����V�P���Lկ�0e�YK�9��qO_L���p��Tu��/8�ˊ��Z��]��A�@(�^�1���s�z��'�l��x�}u��A���<�� m������j��1õ��B��iB��	�A&q��6�t���+�cQ"M	��յN�I/&�'9�˹��Vv�t�R��FAD�/��"������N��+�',��Z.����xT�;(a��C��?����Drɴ��J@a��m�e��h?-����b	���M8=�^����=�ӽ�b/��Y:#�3���rp`��$G7��0_��s�N���vo���B��
]\�R�	�e�1cٝ)z)A���۹����E;DO�V$���t+˾C��@;�sA����.���8yQ\��Gwz�O/9s>u��ř����e�5o��e=���qפkx�t������]�o�O��V��f(�\z/�x�@P�p8��R��fU�j�nL�`v\�\fM����qY�cGr�?�������@�W����:��7[�zȏ����{�N�ND�v�bKT�
{���=��s,�{B-#+�Vx�Z�%��/�(?��9&s4]���5���3\>�P(y
�6*���+����&�sN}wT�$�8���/Aa�ԥ5i[����x@�� �`��������4�nc��,��R���1��q��a��­��[C���	�~n���7a�F��G�S̻1[�#ݹ rŀ�}�uNʂj*�6I�VU˕��UP�����h�1G�2�Rs���Ծ�y[�J�梵3d������A���i(Β�����~\@?�,�8�(ݙ"�i��ݤ�܇^��g�ms*$��ESפ�#-
!���U	�����lQ�̵��K�1u)�ױ~Q ���16������	���8@qY�&C��.:!�6��;c0߷s� ��g��"HSK�P
��10ڂ�|���}��([��`�d>�*��I6�c)<���H[Y�ғ���,~ �lvЧ%	Y�m�[��>+�8U�t�@�e@��v�AB�a������m����p��_ \�**�>j۪��q�E'|���s��}��)��Һ���w,���n�b*� M���1?VPg�>V{���M�|j�:`�@�������x��Ox6���Q���s5��I�a��P��'��C��ݽ��(��/(���Y�<x�̶H|�d��kѺ>�Y�G`���*"�r��l��$-.���A@<��E��u�#�n�����,�=�bB�B��^ͧځ[�<C��^� ��|�C$S+��G���.Ԟ�*��� AP�	�oe���W�\t ��i����� �D=CZ7��<���?��1����m!�����;ZЮ��|�-����;����ٱ��rO"���_�yF�
�`��!�;��U��X���t��(�JW9�~�#&�M���j�n �I=�x)��s�Y��rvHYF|>zBf�؉P�":�m��'(����n�?0 �捻Dr��Ox@{٭�Qh�BU��_FQ��(p��
�zk6=U�E��+��2p����v�)��Y��4`�n}��Ƕ��.E�Tes��q�e� p3I�k	Y�պ��ľ̫�}�Q�@�i���u��<��mЭ�6�e@x~_�"^X��$Ԥ����txY��&��_�/薳�q�1:z�3#9�Sd��V������#�����m8./����V+}����� ��jm�*~Ԉ`*P�,��\aK ������=}�������1�c,��s��E��J��3�2doR0�e��&��}
�)@h��}�G,;�`�͉BJ�Q��ib�]M%�%ᖝ�$�3���0f����9��.����l�O�u+6��,w\μ���� j";+k�Q@��7�HDi;w��d�N�Ž�͊�BX���+z���I��Ӎ�R��2��q�:�r��Ť ꛕ�4�J�\Dt��>w&�����Q�)�,m�k�b��	�KM�PA9A����C�T}�v�٥M���dҊ-"�Ҧ�^���o"�.��Jf���Q�^#��B6��&���(t�f�4��g~yŪ�Y5����A�Epq�3���Ĕ'�Д��*�AT:Vb��|���-%�uw�e�I��UU<��2Pl�SF�׋���t���ޝCɶ]+�7���Ld=>e�_�T{�+�F^Tx'M����DE�o�-l���P�G>���Ѐ]
�?�8a\I��$��B�Aِ�"�n��P�j�����Oy��eDH��t�k#�AX_�&��O�-���T`g��JK�7J��"�Ÿ�(64U��]'�YP��D���я���rZ~�xy���uu$|�2���d~���a�sa�w/���������&���5#k��'+��}PkH,h�d��v���Tϴz��Z��G�_ZN�ad$	c���Tx�4�nʤ��6�P�����ʞ���|�uxP�[�+l��VF�߃)��k�~1s��Q��"���c&�,�Ƶ�ͦ�X���ϠoC��l�I�v�$Fc�I��2!cY����RI����-䋴X�Za+K�k��Z��\�=�Y����n4a��gT���SQM����܁G�"�]������ ��wl�q-��/\y�u��f�ň7'�
�l6:�9��#�!X�Ě��b�����F����w�:N[h�[�n���=��C1;����M9"〧����;/Quu������� ��N�ۖ^$b����|7���V�Â��a��s�.X[�H��M�K/�evTv>�U۟��gSǄ�E�|���Hr2���}U{9��y,{�hh����y� h9��&5�Pg��X�s2� �b��ͼ�tzer��;�4O�+NfpE/�ݔ��(BW��r���9����(�oB6������픴Lq�K���xRtJ�?K((2�~^>��npM��Y��#�)a��ݡ"�#�|�a�*�*�j���[e�G(>�D/��(�|y�W^ x�m#�]���h��0T[fLL�j�~Ԅ�jo�u��9���p���r~��So��}�'�ť5^LP�1��
IJ�p�C2�����IJWC&� ���/��\���=%ݰ�){�����{8�ގIR�v
�Hp*Mi֪�X;����SAe���x$��V+<�$���s��\~�z�}x_a{�x{���#2'ͳRl"�/=?�z`��V��s����8�>�ȷ��k��*98��е��zy�i��S�h�4�?_�\;���Yմ%�V%��b?�����ܕɪq�ꑝLO�t���RT�^d.��p�*�> '����'b�CU/$mް�Q�ql�[�3@��pu��ToV�@���Wz$�jIgg.��]bT��$%
�?�H��4(eh��Խd�,�m��cn��B��
�b�9�uLT3��	yX��a�*O��;۬&����Ⱥ�6Kо�S��`�\�˙o�
��Z�d���%�����隲��/�@,���z��҈��I��cW��f�HЈc���h�|���Z#��Rt�Kj��N�\%�����n{(�ډ<��3�r��AI��֞��C����Gz�.Zm���J\i/��I��)�k|�c����l3	]݄K����'�q#��+��?_v}c�1N(��ߡ��~5�(5�T�Ӥ�O�!��n���0{HMWǥ<�����e��ؘ298���i���|IT�VDb�*y�>w����$�Om�~W�z�n�W(���r�
�z��Kȯ���'�q?Z�X���U/7���3c�n���e�����հ���e��Ym����� DQ� &5��}z)t�ȩԻK����k<�q<�2�1���<79��������8��в��u�F�'Z{r��(ഏ�,5O�o�ܙ�v�ʨ���Sn)ړ	h:ͽRj����D��j<s���Y�H�5R��z=�B���㼌��a�}���UZ�6�@d5�b��	��sV��5�n��7n�:�m��!�'u�	l��1*�Pte�
(���l��U��<$u�{�<l��F@�O���Wyl�@�+,�)����a�
e��k���O�X3��J{n6�Z���G�6o\�]ʚ>��R�,�g.����{Y��ma
/0���U�υWcnI�*%\��W�+�V�`õ�x�����b"�r�=�\����Kmk�)3��g3���	Y{�D�}<�76+7Ŭ柕� o�|feQFW�C�:?��\lS������[7tُ`@?����چ���� }zY��E=	)?YQQ��-ח�q��syBk�S�3Q�0�w����`�ӷ��FI�e�c�B�g�Y���_���x��l� ������l�MҦd� v��q�P�>@_�����^ZiE>�)>���K=��*�ڍI�t/��.%S�B@�����T ��/��GJ�{�fm^ͥy8��ro�Vö�ϿNo����i���ѓ׹F4�6�>jY�::�zֈ�K8�Ϩ]U5�SX��k�<����)�Q_���ߙ�%���sY���}�Q��*��4f�d�Q��*VE�z�5�
xI##:@�t�}��+�{�;��$Mr�J�������/�\��1x��U1y(¦}]ĤwD~���C���ڣ�1��H{�g�d��4=�Qa���M��QZ���ը��fGR�}�\��8Ғ�q��}�4;l��/LoF#�T��7����֍1�ޣ���'-�xT�C��h*��-'�I��M�ڈ�s��/�_�{�����G��L��z�����,�+����F*�޳V�����>S���D�Rg����;�m�.V<�����3�t�`#����N������M1��nܩ�7��u&�]�{جʦXO�k�௛:Rg�L2�4�Z��O�TS���q֟[� ���]�h���uj����X|��Vmwa�O��D�����K6}���n�Z��Oe��b�u��2��A�:vq��L�J�� C"<��Z��������������;��X���H���[���jB?�ݧ�#��Lr
���-T:�+�D֗��@�E�ѣģ�|Qgp=��F�uK�ܫN���Q��� B���Ƽe{\[7ҵ��H���n5֎6�~�b�.bצ�!�P�	�	G���k�눸������J�|������^B�^�Y�n����5��f]$g�(M,���D�h�t`&ȍ�f�j�7���xYg]�22X_7�����=��f��7*qKn�ֱhUr�Y�}$U��G�e��_~�T�1�;��j&�>��!��I�.�*۬�=��(��0T�	�GU�Weh�7bTQ=5�8�n��މh�\�_����+D��YZ�wr��V1Mw^im�G��@S�ɚ��� �w\E���Y�wStH���n�
H����v�.�ѥ�n�]Ux��D^����ї��ox�%��!�����NKx�#��:LۧYf<�0�W�z�4	ռ\agM�*�L��2�^caJˊ�:������Z�&���DS�zu`;%4��P���f�e�`�c�wH}�*6@v;���9_�ġ%�]���gƷF���S�T��0��o����� =^=�
���"�����P8� �ױ+^���#�3*d��T`� A���F�>�o�{�҅W=���ʾ�3�yq�z\�S�Ѩt����):/���G�*����fZ�5q^�3���XRg��X?��p�O����7p*�̄\���-��d[�P	M(�vQ���nS8�Z���j� 4!�f���&N!���[>��^������c���
��Er����ֻ����۠����q�c�]G�1}WUv仓!TE��d�*u��㴧����ag�1�Qz���,���R��yI�u�(֫�^�6_kk���	h<�"��Dk�y���'�ߋ�n�)�k�K�ngX,�h�{�]5Q{�q%��:�Dв��^ndH�P�m�R��
�>lB�D"�tf�����^O3�e�z�stX�g%����u�	��<�W<��m�Y� CDhkX�� ���fß�| An�G
�H��`�h"���L,���;/sC����HL��/�2mnM�� ��G2y�d�of��;���>$�����m=SfM;��&��n;	�,ů�)�Nl�]��3잡�.[;;˦��Ť��Φ=w�^��i^���`�#I������X$���}���L���l��4
��~Ti0�l8 z�Qٚ�(�~�y��H�`i2�>a�S��U.+׸��L��TO��<��u�@����#	�m�s��ӆ�u��*���~��fj�6���>�H+��m�8�B�������l==F���t��'Y����eo���|��$��tT
n���W�k#e��ND�\nB��.�l�,���=K?����p�|[��5��O �x5�L��z�L��Z˹H������ׁ�3�F�Q�Mr���4�4���2k���m)��4e0�$KufN���'W������L��3��̡���i��t��nQ�eJ-�X*\p.22�	`^c�9ν�z,p���ş Ɉn�}# 9|z!D�!J��W+�g(̏���\w��>�����	�O1���.��p���׹��\�h�(6�3��d'�jMk�XC�ݺKc�E���$K8s�1����m0�# �
�Cln�#z��gI@�gAЅ�t���:�g0��Z�2���	�1�6/L��%���I�(.-�}�g�
�)ޔ��}��_���OrV�^���xK(��Fe���^��"6�w9=��1�k�k/s�bQ�1L1ԃ<�)�N������uac?�{kQ���>��
@������R��m+q��j0ߕԓ���	&�Л�軣����b[`�����\�:��s	��G
�� q��H����r4K�;@��]	�D�Ӹ��$�����?�	W.@���)������%Eg��G&�Z�ɫv!%�h~�=p���~xjX��(�߲^0k����W��/	��kмj��P�
ʑ��Sv	�E��1~��R�)+L�
Y�� �P��E������=���WH�zq��{�3:k#� 
<.���?O��H�v���܍�M"r�I�c(��A�5�Ŕ����،�z٣�B5��~��tI��t��X�}�|N7pf���M�ڷ<fțP^�̙\}&�"׏L�p5
x�R�1yQBxV���v�T�%+�������j�n�	��E����#�}�z�-��S��G�=qN���P��76��2y�ɚ�����pQ�XW���4 ȤhS2P��+ZK��s؝ڛ��o�'���g����l~�`�f8)���>��z�����V��������?O��4��o��A�ΐ��&�d������^$�0��ٍ�47.V����9��B��OKH��<*S�����Gy�VJ��Eu8������\����)���kYp�<�l������'��|ݻ�NA~�ֿidC�量s�Tiy�E��r��x�?>W�F����N6a^����}̶Kn��
��-�����>��ݑ�O���ܡ~��3� �(��p85C���pR�n�{D*�Y�`e���zb�1�L���a�Z&�AE|�/Q�%н��]�d'�� �Vx���X����9ݵ/��t���n}"���%c�^�����u#}tD����@OK�IT���͛S�&��#7E�bή��>����գ�$?�o.��Y����DYP1Ёt��#��d �	�F�7�o�vؙ�s�5DZ��[ �w/�E�j�A�y����xR˚���cGe�����rO�I��d���r`�#��7�<Ʀ*Rv-:vE�ُ���?[��N�l�`0��_�����/�����4`0�Rp��3T�z*[�'�L�:��{e�]���z�	��*���I����ފ�j7b��~�_	���8�)��PV�z����D��8����Wdg1|�z� �(�߂]uB�p�:�%��dS8���Q�B?WE9Tt��̀	�ǋ�v��7��,Ö���ip@���ڷ��U�s�}sk���c���;���r�>l ʾ�����K2����"\ف�{>�!3 E���o�.����7��D��vv;��Zu�b�&(��_��eD�>2�H�TA�E#��s�"FhAb@j��%Bm�@�Yz��X��'hN2>��������M]����>�T����.��ʂ�`���<!`B�ju��`5r���`"��$	˔����T�F@�m�\�(k|����;c�XS�D*�}{�!ODC!�x1W`G����a�DG�z��B0�;�]�!� �q�F����?�8K�I��0͠����0�C�0\{�>�'@\�Cȕ��P?z]�*�1���e��C>@2e_���(U$���#S<0N,�t��i�;������'z��'�]�cDm
D��#+R���_Պ�����a^�����J9�
S��%t�p�������9�{�F�N�ǂ��;=�?����_E����g�Z=��;��4�2 ��)��\~����"36�(��C� G�)��T�pN�s��*?O�͂�rd�Л�_&Ϣ�{���vX�v@�;Iϻ�^��tP�����p�?�CG������+�D���o�s~����~ߩ�Y0�4��  Kn	�T ~} T��a��u��J��}Wn���NRVՓ�v��#]��9ʂd]�,Z���̭L Ț ������E��,�/�DM�/}j��HI�O1��س��m����N+?v˶	o�LQ��6�W��@\e�p��uZ2+7�&�����~!OV3�\�Q�c�0۴9����wN]C=��%2�N�b�|��ׂx;����t�E��4L�+��j�d6�YO+n�YUMP���ɜdD�=`` TΙ$(I D�5��^8њR���d�e�ɰ�}v߸п`Q��?��{t�LF�/��k5�Y�#b������&� �iw
:S���\�Q�vQ�a�(��Ͻ.�%�X�z\]��J�K4��}��<�ư*9��isx����?{�㕙* �(��z�׸��Us��:^��]V3�M�߼?�g�皖���rS���jjS�s�g$�e_2'o�G$�����I�w^��'Ӻoh�"��^��W0��rK##��9;y����܅,I� E�ӴMa�sv�!��?�t��� jG�7ښvD��΅�����t����s¼�0�������f�t�7��(}8�"�>�����7��fTP�Y���ٲ����A�T�t�]۪�pq�఑$JF@�@m�M����]��P�7��}���˽S��@O�!�ҵ��n�׹̈́K��X&)G�m?a�S�U#ah%��	��(��+������Gyw4�L7�E�;�r�\1W�}������Rԉ؋����R͚C}Ύ<���:<�����q�\����	�d
+I�~y�<xxQc�F�&	1j�6J¾�8���,r�z�]�U\Уv��.<�M�]���6�����I��B0�a,�[-�����C�o�0�qcè�����t���m��y��`r����l;[��j�7����_�:�����°ԝh��l�k�^;�� c�eIv��9�~}x=a�{R!w&��ݒ��b��v��gO�����\��:ټ�?�[Zڱ�i�	$H����;�\3G�s�k��"h��]3�oz�&@�NV�	B(����s8�WuM���؀zw��(eJ?����,͎ø�o�����1/�ʙNك���A�]>?��bby�H�������OYjŝ�.~M($k*���AD����9.Mn�w��sۭ;��WJ�u3�j�o���� �8]�Z��Ͳ�`�:��� �1H~kȃ���h�g~ã �m{�xJ�}���f�;_^ܽ��<k��>m�&p�h�������1SEi.Jƚ� |N��0� �#�i���_e����{+/"4jS��O;>��g����rAlP������/>àÛ�Rʓ�`��r=����*�U���G4��_fx�"�Ǳ\�X�A�9۱n�5���1��kЎ��y�-��9�1t��&�=�����hN;�}�.~7o�qU�+��照E&�V8W;Ͻ>{PB��ދ�z&'�������	���t���LgO
�,�9?{����@��`�7��������!���[�ʔ��H-20f#!)�99R�4]���IQ�T��f?� �o�3��>�%X0{�}�R�2�GK�W�5�l`o�AK�4H/����dwh�>-�)��o�C��.�r�C�f�����^�b��,9Gc{,^�9���9�u3����o���&�����j������-�T����،�=���t��������`�T����=q�����bff^���@�ԧ�m������_�ܱĂ���H���vr������=�q	7�Rg����_I�/-����|؛�>uɯ��BQ�o����Eþ�e�����A�!�;<�uz*}�wa�N�����&wr��?ȟи^�v��`��ԺP��͂�OB.�,r���	�߲���q��9�?;�Hs1��s��#�U�Ӌ��*��2�o
�n綱� �7g��J�-��u@M�q����"��ׄ�v����Ղ���vW�T�$������S���N�:~k�m��Tr��X?M��nU����a(��̅��o��i@��[����pj�rNpX��W��?�h�2�2-���`�W��/��*����؜Ps
�8 �� @��ݙ_�c���5�FL����;qA>� �k<~�Y屼�G���ōv�Y�7\/䃧�F�J�8O��.�Ҭ�w�;^���ӥ���64_�����
�Ƨ�g�l�N�]9�z�N$Pn�v6 ��ƤK�@���PZ�N����fM�*!��}]��`v����

 �)!���2CJ�����L���Ӭ�>��뭠7���;����@��egXa�3��ay4�w��)��/|)u�4��3��]`c4��<Iٰ|ԩ��T��Z�#�l���q���^�������<r�3{���;"��
Mw�����k���L�j{���i1ڕC�ch�3J6[�#Y�
�o�i�f�u�Z-�@���|�.�g2��L>�	����ʰX������HreA_�pw��[&�����_�{�Wq��pL{��U�w"��RMk����2�zœN<��>�4,M�z�B���~"�_�z|
j�l�T��Q����?{4�����~N�_�ƢE�v��H���ϩ�#��GO��M�/�֑�k�.H�s�>\s5��I�&ڇX�̒��g�0���u]^;��d:�����S�K@�#L�{�od�F�,H���c�\1sZ)5���u}�{B����L�5�?�T#^�:G�-z�u=�ь�FG�C����s�u��j샱�'��|��{���C���|���<$11��];����#Ъ��]4;�V}s|�f#���|НS��� ��m�J(���t55��E��8���K�=�)N&�}���U(�ׯ���w��(����;�%�RWu��J�Ś�I��~��KA��;OV�@�~>���TI9�cz ��*@���򈌴(��	������{��Ps%�n�E��轶g�;*$P��U9��5���_����wU������޲��*�w߬�P�D"��f��"��\v���i��T�ſ�D����'л�?�?�c����������!��*�r��Z۶�+����8�W��N4K����0��P�=A�Id$u�ߪ�-�S�y���m[�aT�����Kw��x_�ȷ��j�������hg����=���������7�0�4�1����@48�Iix��<$���1I��gb`/�V��R�l%��'�H%F���m��=����[��=N�\|��(��	/K���J��γkpۆ��ew���&��r�1�Z2���@`������lbj��/v>��y\m�@�J�0�,!�r*o��)<���QqaaÝ@	r_˦K�d���$�����k��m�=7�8�a��.ľ��S/�F+d�d��]���_���9K�9�ڼ�KO��D��sh�����=}|e[�K9{U��햲>���v���8�O�ʥl�U[�Hx���$��Y�/\��Y�$N����F�	}}P�!���==2�:h~]����y��cQU�ք+�5����LE礮ŭ���
�&3���O�R��u���`HUE����;��:(2S0���1�|�Z�RTW�[8{0M*���+Aj?���!nm�4��&��9���CO�ZF�v���|��.�^�kz=����V�ϰi��=�։R7�|�!hR�� �Ra,�7��&՞Q˺��.��#�vg}����2��B"4C��/�̵4�}�QֻXل��%oj�@�������h'$ЪX:p�¸�wh��	���t�'/e.83}���<.�;���8�U�z�������"���==���ӳ�?Β�:+���=u���oS/������U-���?ǳ{�)9����:}VL5�)���^��.��Y2ri�g1~��em/�{�ȅ }ȉ\�����ޤ����� ]g[�M��޹ժ��q��$�)]����(������)���0��j֧�Q~֟Y����A�yוGEwThe1/�67z�ظ�H�J(�''H��t~Ş*���Ҹ�ϰL�̐���!U��"�Y��f���g -����2���j̞�(�p��0��]���v�z؏X\���̫�=.�jk?��[W�V��o��C})M2_x٘��-����|1�<��JU��''�y����h�P�W�#��������bvM��e�����ְ��2~��N� ��M��F��ͩt����ʼ���F���U��y�\Xp	�Q��uչ�0Z�*�nԔ��;�!�k_��CN��x�E����PM���<��i�AՓ�"
����E����������^��7-�e��ƙd9ʇ*��x��JcJs�>�ԕ��M=�EC?x�#\I�g��3U�{7&��f=�Vwh� �l\l�h��t��+��
8��l�e��h&���7�<���)�'�Kf	����ːDz�r-m�C*d�dl�ou���"(�bV��_���d�#��a�4�`��O��%�lӑ�:
)����X�B*���������RN��
��sƁ��� x�)�+�����.G;�G���q�_����F�(���G�~��>�~_&�6��0`��(�[�\�N݂]\����t�?����s7^���//��s2�PK3��� ����C�FC���K+]�)��GCi�H��tG
���&O�ݕ�bֽ�:^��6�R����$�Ԇ�Ig�g���Q�ˣ�j�W�OX��W<�����DX|�����Uu���qu�	k�Je�Xpӕ9��)�d8
�Q�a�9"=g&���A4��wL�|���g!W�<�fJ����oh@|��|��N�`w�;{�>�r-W��nN�	�M"�}i67���#Uvß���+����eI�~�]�3}�eC �ؤ�qc5�
Z�:�z@��5(.�Ƥ}k�Zs����J�?1�7k����<�����xf�	����^���$U��.�Ս�7���7��q�gV�g����t��Mgߛz���j����Q�?:��������;l���0�l)�J@�@X��'��jwx��پ1`��p����~|�<�	>R-��鞬G�M$�_x�i휱g�i�
�7$ cE��ɸ~�O�T�L�I���o_����´�nI�y�/$J�L��ȆA����2�׿�F�GF�=�I	��a�_r˟ ��P��j��3��q�iL�N�����$��/r�J�o|���~��bMuuC��E���%�[�*R�{�����ĭ����c���όI����K ����u:�45��i㫴x���CM����8V/�,1 F(sa����j}W�I�{ZH@ڃ�NL��zxA'9��p���PJ���`|ĩ�֒�h���CO����t
ujL��Y�7�a����6�����w�o�x�3R��J;���t��h E׸���z���7�KX'�x��ڢ�ULW������ipw���x�M����^]��;:E1�b3�6��t�'�OB[�0B_�i�6���,���Y.L��y�ܙ�F�ouZw��O,3$m�r�}��6�>Cx#��t��8�����QM/_ߨ�c��X�
�DzWi
�;��^#��HWz�{�� ��.%AZ(!�����9�G|����u׻�k=�יٳg�ޟ�e&|gB�/�!�>��	[�^l�I��۔��<$� ��rŒǅx
-V�-��T����T��h9�	��oXi�&��I"���yEH�;~�.k��b��MԊ.l��d���u]���m
��3�����8'	�Z�s^eh�����<9�hW�!j�S�w+GǪm����o���%��#*��x�������i�]Sr�ytfh<Y]�4��i?O�R�/h�7�$]��ث�f��\W�=?.-3Z�X��e�.5���'��8�o���7�zj�3_��g�E-S�a:k;�o�3]�Q�j�����������&�y�b�kJ�:%�h�R>��9�!j�+���� r�)��(�8}�S�۸np	�}-�hI� RT�L� ���<���fH��n����``դ�+�r��E1l<��
B���LrB����G��X�c�[Hd��<6�� �/o�M�R7.u�����qt�i��ǰs�3��\��h�#��ʇ�]�k��|~;�L��y`�0'�D#�L��J�""*��#r��6)�^!k
�����`O�Y�0�m�[����Z	>'�g���])7)I��\��6��*��8jO�SjB�6�ȨUW�m���Z�=��6-g��X4OK��K!i��@mx��=��:@����"r��CE��"��i23n��FƬH�S�U�Ca���m���Nc9R�i��,2�Rk�4>�y&���H��^�OR��cl;���*Z
��Y���\��&7�X�s�@��w���Yw�~ W�Wǵ:���E�B2�s������m��#��jz�}���rV)�|+I�յ�y� ���7&06�5}O�U��/�a�+�~�b�m_ �f'(��޵_i�OR\n�@`K��p����>�ACf�d�<�j�wgC�_���B�)��6�ͯ�ne N��_�FA�sRG�{ô��� >Qį����U��:s�zOp����551y����8́�����G�������.�k�5o&���(�Ɖ&dd���F+�q�=�Y�"L_�G"2,�T�嚡�'��ܵ���)p�`��p*o�C�EB|s>>���!}t�挿����qZ �\���mK�W�G)��|s�Ɨ����s��k��s_���d��#�B7�1�
lBR�EH�u
�|���ǝ�Qe���%�Ñ�u���J��%͸�4��O������~�"�͢����#0�OHK�ǃā�8�ǀ^�B!}S��F����Ȭ݈��j�ykG{�A�P㞣x
�o�USu�Q�[��ټ��!�
e�T7f�<bM�īvk��ZȦ׀�Ɇ�j�$2��N��&��ϛTCۻ��o�&�k/���u6���[,���6!�2BjK���x@�轅+�,;�2ʻ�n���úL��ب���:O�Yq���5��+]}�0�b>M�[��V5*VRɄ/���ARՈ��o	��<�v:|���`ϰ^Z�ƹ�I�C���ܝ�:�TY�$t�Qr)��}�jM��CTS�k���v�1�諸�[�b��nv�;VQ�resK]�\n�dG����'p�b�V�L����k��m��_���[n]4Wh�gGi8�"RW�h�n�ʷ�!���Ş�$�3�n�w�-��"'��4��o�	�YWB�H��#�3h�D��_�mA.���9̳%��q�Cb���{����Xrz<B��f!��E��[+tX�z�(P�rZ�`��z��*68���E�m�NY&����n��<a}�(�j��Od]KA�vN�>�e���+]�
s���'*vP+�>	�-�6
�[d[��Yj��oh�*�кT�:z;�38߲� ���ƒ�8k�vW�7g��[�7B%�c-���M�M,�*�q�L��.$��$�w�?���=a�Q���5)�$�
ۋҰڞ�}��s���lU���^Dg)Ќt�q���[��������)�&�>��K���6��FrY�`{|QU����=�20
 �*6>��$�O0=�U�Mbّ��L1%ios�<p��l���ot6�m���oI��V3b�xҠ���W��Ob����A未c�[��zq��8$�����:Ӭ��\�o��Bܠ�z'|���I��zẶ��[��5D�k��+��
�J�'W4�����yߚjYE�l�%6΂��{#��+�_#�{�?�9���X ��}�U���n>g��͕�x��C���Z�~�9��ۮ������DX;h7��wH���~�@@��d:t���@��%�P���i�Z�HLLY<su����u	�⮦1���}qa<o�x�9�e�?n_�|�RQ�
�gT�>�g9z����j)@m�T�V�]�l/&�~�r.�*�A�{#w�dլ|�:D��+��T\}!��³���#j��� `��:�$k�ڎ��>0$�<@s�[�9}q
�K5M��$�y���"�'�k�Z���E��M��|c��:��+w�e�@�a|�;l���V擖�:]X�b>TVw/�2{��)��5ta��U����.�k�3��w<���ٓ�ҜD�1$��σVk���k����-�{������#h��6�ŝ��LqVuSU�`kN{�嚰_�M�.��}�@}��ul���Li�S��g���5]�+�-��`YTu��x2.��e�̐hY2�~�=�j(���UU-�7�&|����Z�"[�%���dt��W%Me$��ɒg>|��U}Q���h��{�=�4G_��x%�1�w�^��R�Wy�[�̩h�h��B�[�B�U�r���Dҝ͞��V��-0"(vߍ��X|�����*���*�l�DS���d��Ed�L�[�~G;�f�Z-�ж�%�Ȁ�|�>�~�@��Lh彈��6z��Ͻ&	e��J� LOot�:x��Zg�Ϟ#��(#���.�Y�L[� kC�ի�.������|�륟���a5m^�:V��Q�T�c. ���X�	�BϹȂ�fe����99
/���YZ�h�c���Щ��A�ac�fӢ���ojA�_�b͏��������ߞ_ ��z��I���:/ r}�,��C "l!w,d�{q|��Ǟ�������sVα�m>�Z�D[�N�85�
�m<Q����)w�������C^EnQ�S�w2��X�D+��J��0�Ub� ���Ė�S��r!-f�X:m|×/��R9���7ƽ�4u���]�&�/i���Ѵ�>�`�rX��,�,����q�ߏ�����jk�4�������$S�t�Œ�����o@$�q-��L�`6�L��Aig���gc�ᶂ��p9f���:�����F�i��}|�.��E��+�ɴ��[}�!�377!V�W��v� ����(���fūj1��i!S��w�x�=x<)���!5����~U���)Db�[f�:S�i�4�+Ͱep[5MS-[f;�/-�4�S�mX�g���e�8��E�nIV�߶��<�IR�D�+��s�
H��ZU0���Q�㙹��%*�D�r����-���G���w�����׊h����a��-R�U ^z/�_-�]y�e�8;�M���+_S7B�4�
���Ro�y�m�+?	����\�ݫD*�_��&���NI)�;t��&yñ][+�"թ�!y��˙�z�Ֆ$YC���0�e��[|ح1ʽ�y��OM�zܭ��|q����VΦ{U�Ѻ�z��֘��XS��y�"|��;�i�x c&3�ڷ��k �Oi��[ׯ�6�m3=?�U4�ݴu��x��#1�x()=ׅ7��'��B� ���Y��idr`�X�oH����5�2��=K�hla�h�l��MY�^��$�N������Y����*�� �R+����-;��ؕ����kƱ��[9���{o�XV(����P0O~����NV c����r��S�E��"�6���@����w��Z݁�#"]�b���)�(RazG-�UC��gp]�9%�dw�r^)6tt��pҷ� �7��uX��g)k�5��q�x��G�
���6����^K���x��0�c�sQ�&�H����a'�7{R;���l?��X/����
Q�^*ik�����8a^s<e�" ��N��-�9�t��u��!P-�����'�CAէ�W&�r�+��f��]�߇%&a�k>���>֯�����JW���U��Io�� ��^�������޺�ni�o��t�_T�u7-����C�$�H�l�7w`�k����Q0 S�[�f��~��I�\��Q��'�6���L[͕6eE���*�#��	Q���3�R?ې�Q��"4[�3����ʘ�Z���eM"��\����.�4�\E��s;Q�i~�%X��X��@�G��?�9e#�~ �N�DV����X��&;a���L�)��6� b���w�9�����:��>z��w��7���C�5�&_@�	iI۪�|���F=��lG�2R޾�wyJˑ�{{�̱O�_U�S$z�3�O�qЫ���{���E*#1�x���P$G����GƄ� 5�M�'�<��|����9�SLf)�Dn.@K�׬�D7o�Љ_��6`6�^w Չ�� �2�+� �D4��(�^�m������@�᯼E�'��C�șq��d�Ze����D��]�.�+����:�t��ʐ�5�>�M�w;+'v�pX�<9O�������r-nst�o�Ho�P�����ֿ�<�H�LW��Z�eN2��4���O����ؕ?�{?�id���;�9t5|�0��M����'!�O~���ᰣ�	����E�>����)c
KV�z=��v�cv4Qm�]�%l{_�/���J�z�DԲ%�������T:�G�� ǂ��-�k�=p
�h*_.cr)���b���n��B�����M����ŝ�@7wT�
�*�u}��ļ�>�Hnd�m-��t�S˔`��mX���?'[ǭA�64�3Q�E��u8Έ~t5xխk-h�3��	���f>�9�r��i���t�m�W��x(��;N��&���C�ig�L�K�yeMHJ�7+<��T�I�������U���o�,���[U���@l{�zh_+��~��y\T{�Z|
AA��S$:w��	!�YUa�|�u��C�^U�Ms�����Z�Pqc9c��V�/�a)�
�~�F<|'�6%�jk�)��@��v��x����6�E��EK��+�rx��u|PH�	Qq򉶵�{�T����O�ԽOڵ\pL�Ś�%��S}��pKqE����'	U��8VP�s0��\:�T��5�(<��'�K�Ι���5.�������"��U\��H��"N>X2��f�p
[�e9� OF��4�(ܴ��ͼ���)��t2a���(��R]��*�
�2y B�0�,�
�I/�{_/��bsw�y���??~�U[a%�3`+��կ�DU��ǧ����>��1Q\��
�l�����<#u桅'�G��3�������@��:�[��Q���a��N��м}�Ĺ�*���&W,���.�8Җ|�t����%U�Bk;ij��gpM�̅�v!)�\o�g*���bm#I����a������P�!;�X��Qvn3OU�L<;���tENe�[�@fv�p �%��s=yd��ѥ�~��]�]ҹ��N��k<YZ��Tl��c1���1e���\@YL�Pop�R �[� *�솆C�XS"��R�O'� +?/��$���U����N�z詡����-�Ƀ�-������y�z ��`o w�ne����~s�>���2��Д����R��+K�M��]��tų�Ӽ�%(ķ,a���5)n>5ޣˡM���	>��4���;��N���R���2��R��&�b`�\� r,s�����e�$��D2�ɑ���jUG���{i���XOmu��[���T܋�3V��%_ҝJ^�:K�2�����ƻٳ�P;\�~ϔG�)�Н �|���R�����m��r��[W꼟�Fi���ɯ�6�|�^�^ee�Ʈ�trL~'�݀���ee؉)e%�X�����u{}N��:�!��l�4��n�c���b�܉m�?��CN֖̂Qq�?��@�^>�f�&�ȃ�[o��M�B��M�"xj�O���l�=�������ǣո��x
�iǩ8��|��s���׶8iw��L|_u\�����c�"��il�1�>?�*5O6O�@�����H%r��M|P�6n;o���-8�BK%_	I=~܋�ۂ@HSVAeU�LV�򛊷�y��t���=ҫ� ;_p^y�T)|Y-ϻ����\4!>��z�B.�|��҅�<3{z��Psv��Y[�Ϗ� �L�6b'b��:ې�싮�,����=���7�$��,'�1w$ׅ����C��6
@�9�J���F%Bt]u�*�+���4�#@��߿t��*0�iZ��!a��I�VjOc�т�qq�K|9��'�Q.4Wڐp�~���D��9�I�)�y��N�
Iic��  �A!��n I�p�`�p��[q��9���6�HV��`�WF|	AVMw��/��H� �QTJ@�˶+�Zt��5�f׾�y����8	;`��H|���a�zk����'ʧ처�S�v �Z?fIﭠ�1��k� �X!��e����^c(D����ߊ�y�E�A������F���)%*J�H~DR����K�I�,ѢU��A��;a���j�]��-� �0��6�%���YEb=xk��5�Bt�h�$��R C9���N�����ҧ���&Egc�)��7�:�(uaU/(=�H)<�ꂊl�\^����L�D��JS�G*!��Թ����6�U��O63T�����R�W��NIt�z�sڱk�`0�-3	 N�1y�S����3�"�꽡Bg�B><4�d{�$	+b�Xez���zԞ$@�	K��2���9�:\d^_�݃"�u,Օ��n�UV��Rd9��s`6w9[�� g�?l���R��c� �h���cB�b�������^��*�q��9N���*vLZ�������e"	�أ��Kޱ��$Ia*g%��.��9���mXj���/�1�j��@p��d�f񑈂�dʗ�X�S:�l�.f�w�e�u2�߾�dr�}�<(��1���k�}��sJ�Xm�̩J�.��`�GGr�ԉ��@����]3��������^LG�e��O�2G�n�"�� �7��aʬ�ry��7�ۼ��}b!�����Ĕ��e7�WW�Uq{�H9)�ޤ����O�b�G�x�T-�gK�'Bh%j�2��>i�����ȴ�cJ�/De0[3���c���p��'����ȳ�N��&���%H�o���3s�u4)9}|�=�*�,qV����߲{�+�[���_�L��XGY����d�m�nz�ƽ��%U��2�Yʹ���c%$��Y"������C�=�`���Hy��*�C���@���s*R��CDÉ���Д4��� ��9|�)��׿'I�.���/�g�}1���������,����j������ ������~������I����w^b�����^����?#���S�Bw`�������86�L�C���0����^���%���|q���9=d�4�+�ލ�l��!��]�dϮ�Y��5�:���-����%@@f[�J��'����@`�Z4o�k8gԋO��>�F��$_Uy��D����L���o�soߤ)Qˍ�1k�T*���Qd~����'��<����c&%>�:�=*�k�-�2[V�z�>�f^���4}'Xh%�3���Ĺg�X��~�~0J��d���po޶�ŉF&)�CZ�&�'H��JP}�<��f�*'ihV�����w���D�2����}����C�AA���Z��U���{�3��߭2f_�N����7P#:\�`�[�Z�ïa�8�}�+� ڟ�*��Y?���pMv_)��2�Gz5Ri6��t���:v1^�^D��lk��Z��$Iվ�WJ�܌�v^K��%li����~\�x㓈�v���(�!�8���w;�E�&�T�������
����Z�+���^��s�c�z�A�Zk���[UM{�����{�a~U}	�g�0|���RH��^��� A�|$�x�*�Aά�����"vW�n}#��r$Q����@v�&�4�[{���Y�غL����M`���Q$�|xq�xR���#l��#J6nf���̪�J����7�V��g{"���@��}�-|*�&	��|�y��
8����s6�����e2%��
����X��C��}�U{�T��
khO��
1���C����9�p��
^����:ع4O(�mJ�A��g���!���{���+�M3��fP�w�&�OG?�|E{Y(B5\m�l[��'��l����Zo�ը��
�����aJâ��K�M&5�-,��H���md���<�j||>"�>_�T�r����~Iq����[�}��Hy�(TM&�`��i��rGn�t����,/2R��!c�V���{��{��۲N�ǈ�@6p��&���z�F߷ �=���!i������S�c�2!��C�%Ȃ��;z�b��c@6X�=�j�ve8����4i�2sF�೩����(��"C�À����a���`�����pn�NV�H�p��C�FDD�33Ծ���h��AO��+��e�&���ѓ�)��|ȉ�B�rOxC?��D�����9@��햎ײ6��c'��y(9�a�v�hV�黎�X4d�j�;�����+�v�T�����8�#Q��d<���õ���-��C��&���cD\D��O2�����+�`��J�VP@�́��Z��!��6�juu���>-GkX.&ᙑ��0�hw�¼TRp��W �W���u{
,>MaB$i�R;2rr�Za岦HUϖ� 6r���-Y�tH�;+�e!�������wH�@��P��|V#kV�ݬrO&1���8�ٺ�Iص��$���?���o�lg�I��D>d"���L����hM�b�(˚{
���ha�\Z4\{�*4�@n����k��i�o.���8	[�t<��q�(C�6"��T[$��$�d�~6<��RL�(��Ob��)��\ �J�]CB9��e���n��,��4Rqp�b����gٿ���T�=C���i��{�l	�Qv?��Ņ�W��r_�C5��;�K��V4���0�ј�[�﷏�=�[�٪�����ǻ�Ʋ�~=y�]�9-]ћ��f��f�i�̺!�	�b�E�����(w햾�w�Oy�_iٵjﾹ;)���}|��8jt�Qvɦ-� �����OD�����gt�m���'�䞻����!'ݭ��ok���W��Z�N��}k�L|k6' ϻ��~�����銿P?v<j�J����?k��vtH���J��x��*D���E��.r_+^�����D���+���$��[f�;SvW����J����t���5�����U.j�	' �nw"6�@�����0�W���,�+>
2��씎E������	���QI���0��>�ik�N,��U#���p��r�p�ũ�V�}����o�������� 'q����,����6�kLW'rx��e�>'Q�u��j�����S֛��������a �7��
�t�Y#>��#�5}Oj!غ����ݨ*�*%8�U@Yp�έ�njg�ԝW���a�q1QG{/�-0'D��������/�������L�/�V7=^�{:��R����v�cJ�h|���\G�,���SSo��*��Y���d}���iX����wT��&�0��M����� ��U���jq�6eA�����|�H���B����� ������!<.���@\�j-$��%�^�9�M᫴/T ���ơ��;�}Z�Eҋ�V�9Mm��և��ߤ������TdDT����i�0��9�(�U���YH\p�f�ïL�<��,�����NU�1�bg�>�!�7�W��8~[��!҅���<o����}O��А�]�������i'����:=2��m�^�=�E���4;��z=W����t}���B��#��%Mb+��k|ޡ���	��@�PuZ�l�ע+Wv�y\�eWf0���:u�i��b*p�}={|2$ry�2_�ʊ��7���5��1��&�ۯ�����uK;���|5�=y��4�5x�B��]T��y�(B~TOA8��6���$N�p�ˬj@ZyvHh��jrM(b���i�>����(���-kr�TŖ�����u��Ğ��*��z}��k�6� ]	K�~Ř��p������=�.O(��~�[��Z�����\Ӣ/́��/�ii��yը����O��%�[A?�H�>��䞿N�%�8&�IW��ү~m�Sǁ/���ܤz��qG�Y�,Y�n��ք�zD�!�����e>+P��vʫ�~�=������T_�e�>��|�wJ�"��z`�T�+�;Ojգk<ޱ&�]o�Ђ싮&Z�2Y����D���)j6��p,*��֏�|(�@���E�?��M_�[ �*\����缋��zE
N6���s)1��6J�6�������rDG,���x��Y�Jջ��iЂ��B�|n�E����2��4,�iN�Ep�݌ii���T1҅T`���]���W *����oUS����ʆ`��<X����3 Xx�b�@�!�7�\����!�!�4��3T��hF�Չ�bx��M�}���i�K��+��
���<i⦛I6NCwz��m�v�F#�R�r��5����y}ҥ���7��N`�*��½���s�O���3Z{7+-��8��ֆ�V��Y��7<�i^��;�4eP�a�hi2�2���ᕧ���~J���<O��%�Q����%M`�ƣ'��9c��)�.Þ��Z�*NÞӒ���g�6D��z殍�:;b3�ӊ������n�e�秫����\N�`�9��������<v7���Ƈ�$~o�y���ޢ�:�0g�y�%0�w�Ea��9�^伛��a,�M���;���P�T�)�3l�%���q�>�S�߽ݱ�������]��'�?�)�g26�7���`���D<+.��ۏ�?��L����)���DN3�����79��<�ʜ��%�pjʤuֵ����	=�n}����M�S>�O5'���k�1v�[Ke�vkS�.�����ݺ�)(,l�1�����h�5',q\�MgX!U@�Ĭ���5(��{m���W����9uSS�A��������k�r	X���A>�<+�U@��tБ��=���̵Y�WB[͛�$<K����EL?ui]̺Ӝr-f����w|��*��>W'V5?>%��c�F����LR�u��4ۍTa;Af���G���*��n:�R¹/�|���8������[`u��$�-���,�������ӞZ�0_���� �RH����sԲ<�<���GaR@��y��+	�Wn�?�ʜ����%h�!��(�l.O~��Z��=�*�DI�]:�S�G�`���Nd��������kVb�&gm� ����'Y=�hO{Ƽ��}���N�X���
�����[�\�����?t}�V�M�0C���o�\'�>�P�?��d�Qʨ����1�y�[�)G���j�n��8jf���z&�Q�ityr#�Ϯ;@��IׇV���\�|ˉ
�|!�$"BWɱ.׆(Y�Y;+/�x������^���z2�U9�V;��m͸ں���Z��+�Y��8��>��-T\^��T��Џ�䝒cq��R��m�\�/�5a[]��m,lEJ��Y�Э�4�9�ǲ���c(����_Y��[�d����B�}v{�x�f��?���Q�������r��FW����䙩��r��`8�礭��kK
=��t'x���-�p���Q'</�+))Io��N���O�b��A/]����j'l>�^s����Jٔ�hy�ONӽ�g����ya�f��A�C����'<�.�� �Eq茈���O�/ӎ���%i���63�����e�c�~}o�>ͩ__���i&F<���W��i�;��ӽ��J�u}�6��Ox�衉L�n}���>Gu��(g�ޝ��[�O�D73�jڇ�����?��L9l`N�~���@�J���Ldtt�#�^)��� ���`ϵ��G����՘A�{~�]i����z{��3ix�U<1ES#{Ү��Օz�E�i$G�׉j��5��ΏlG��� ���QZ���B�]�Q}�~��Դ]4bc��X�s�����JK)X�y�ݑ4ϬfEۈh���Z� k�iJ0��6+J�~��I9�3�1����)������E��(�ds!F���pv�쌘5���^���y˹��4V@��f�b��#\�~mmm�di.��$E��/��;i~dH�'���kЍ�&��K`0��Ȅ��$v`T9������iJ�w���]nz��?�9�iv}�c_D#�#��� �:�����N�>���L��c8���Xdd�ܑe>�<k���MrV������P�;�݇�9z��`�Vs�P*�ƳcQ��=;;޾�5�y�.�;9bؔs�ڵkĦ)^>>#E£iJ���-����BQ)�T��Shcy����]�X�&L8��M����P�@�k�#��������QUMmֳ�d컿�q�<1������5S_jSߍ�_���@��5���1��!�6+�MS^�!�V����f�L$f�/uf��)�n�a��]�_`5ݹ��3�4P���:&s��۞$�#�7;e��t�5��\���gmy5�5k��$Tf"�C�'ݺ/�w�^\�|j����K��5-�*R�@�7ä#n,J�����p�NJ��� (l �!�TU	w�^7�t�KH`��l�%9��_?;#�+ ?6��N��g�Nv����u4����e�d ����uj#t�jCG�l
]hQ�A��陘�\io>0�244�Ƹ�O����t��ׇ�\�Ħ53X���1���dB��8c�O3��,�ç M���K�����0B@�!��R�GA��۪|Ǧ�� ��T��$�۲�w�G&� @Q�m�!D��N�.�y�Λv:���`0M۵��ݑ������@+��6�e�7f�SRRz�R�(�Gp���L䔖���!��e���?��F������FH<�i�|�y��n�%�,/�.�y��1C�-kdj�/x�HR�ABH+q2�;��}]A�f��<�:_���jW�/s 	hӯ�B߾���<ӛ,�ׇ?و>�ݞ@�_E�n���^�1����E4탊t
�O9�`�m�h4xm0n��]q�{�`聑��z穆`��mf8X��w����!t�;ݦk�w5�1?7�K��������"�[�SJuL���#�c4f��C���0W@� u��y�ޞ��Q~%�X9�!�~��+°�gv�k8T��y��<�"�i��xe��z����i~��>)""bfq�������ג$���`������?��������Z�ciP�a�-jj��s����Hg�b�e�8��4�d�FW��ו��Wk
��.N֗���</�{7���B��<�#[��wt���r�4�Hp�~oy��Yb��)\s Ja����a�!��K'�!�F!��ԿkN5��5��f9�~���fW�A�B����;�q��4��#���5�%��y�ɺ���ݼۍ������,.l��m����Gwc.ǜ�>J|� ����̧O�0U=����NN �0ź��Ͱ�wu��n��������i�����\j�+�9?���ܻ��.o�P�>|k��33\�~��S#kQ#���ܝ����@��XǫS��aL�!��g�ai��U4B�	��e�c>l�1|I�N�X����7�1}!�ߩ��s�{�������xえ��ʭ@w��&��-H�w����[I���΁?����.��~���j~9�k�_�\/�:�Fs Q�#{l���3���.����us��=dJ���J��á��GVN�WjD����"��O�?ן
=�ރ�0�a(P
Ŭ�f4�72u��F��4�,s6oJ�(�j�� G\�%աV$5�cI�'�;�� �#��A��i1�[_Hc��G�N�`6�N�W�68���!�� [�q[��Ą[� U0���s�Y﮻3��̑�3^ 7X8�:|bpp0P��� `�����fA̛f��/.��{_G�����:��*ۀRpv������	O/��A"1t�]��JO�ز]��׵�k#�#]�ă��*�@f��� �6�0��U�u�FĕK���~7����y��0`��r�գ�-��uu�&N���l�T���B����>bȄ;����*�s7���s�K-�#�K}H���V3E�B�w�q2�1��o�\��^�4:qFu�R�̐V��iAd2���%�.|p���S��[�}����AT��Lp�]�#!��5*��pM��Xp����#�rt�$���Z5~��>�	w�e���C�B>�(y�i���|�ږ�C��ߵ?y��[�D�`�(5�"��i;ފ��̯�@j6��i��V
��_鵌�Z�o�d�{W�<~���E�#h�l��$�\jTS�8ɥ���Lpв/����s�QGBنPQ�EA��7!�����k�ZD�+B-�f�c`޸��t�"o�T����'T#8>�F�
����W8S�����([U�F 8J������k<�o'�n`�����3��kߍV4B�Y鎬��ݻ�o��A��7��N�T-�F6���g��PB.;�*��J9�+r�/��yF����X��8���zn�T���G<�QA�a���ܩ�a��^��,��
v��/��sFiՇH���s��>�q�'+l�J|�1�d������B�xvv�DyVPa�R�e�0���6m���M]<uȱ4J�c���X���ɽ�eUs�dnGAv����p�� �R����9E��z����fEw�W�@��.�1� !6I��b!�HH�R����5.h��K�0;���1�wO�"À0����N�s&�1��5�F]�Y��Ai,�Xƨ���2�ʉZd�&F;{^���}iuv�{s�3Fri�?r0rf��$H[�0ȌX�D+O�;�B{��#�6[3�x����V:�@�Vz� ��:��X0�r��2��'��
˄*{Њf�x��	O�gb�N���O�t���7^~f��B�|���l��o����D�*�R����l��/�gEWk$��r� t�OL��˭�9����i�w\jN�\ҫPS�4�*��6y�`��CM?ɛi,B%$� ��j���oȥf�@���x3���#�;�Ԝ0�A-�.A'#f�VWW�b+���m& pU)�rt���f�I5�yp�<@r����� P�O[m�un�D��v����$�Ù����v�����*�I���f- H��v�Gieq�(�xfZ�8��ˠE��w?�a��0�������/�������C������xV���X���R)oeH�D���>�7�D�ĿI �f�������B�P�_��kte����
(��M ˰���#<ѵO���Ȉ)
~ix��7�]�]��a=�p��������ֶ8�wx��r���QGy���/S��	eh���TR�_���,��@��@�u��31a��~Y}���'p�w�^�����`C3ޕ�~gL�swt�%5�H3gۦ"��2����܎G��.�|��?�.��`�/�A,I[�z�4��eʯ1�+�s����8WY�Ɵ���IE������	�i��+�R��p�6y���N�Ǌ97�Šo9����!<I4bsrA��+h]k:
��5K��J�L�S����:�y|�PF���O?�mɓ�X����_�'���yY�/�mG*� ���$�d�T�p��d4��?(�%�nx,��)�+)� �o�G��d�F�E����;��[�*#���s�L�~.�%���lu}eBr3�>�t�n�h�z�pt��Ȧb�vK8N�`�2<��F��3���eƺK�d�te����6?�س����{�G�7��e i��x�r��椄��Q��$(��P�}>IS���%�'����� 	A��Ί'R�q��3G�`϶5N�bHT"�	��PWJ��A�/�RM��G����EN������
ZX�X�^�i�_ڒ��`�s�\U� ��Dg����B���3�&��&�0�+c�v��\BQ�v�`|���Y3�_�4�ܴ:�s��]��/��iǀ���|^瀚���)p3�!����_�T����_��_2Pל��z�+��?A�_�����s���1j@��?~�e}!j�B�GG��$��?Ww�O���i����E:������6}�:�ԔRO�޺����ڰY$Q�8W͘)���J;s��٢��SCr��z�h*G��@��������V����{q�j�.,��ڤ��࠺G*�j���[�>��ͭ,�V��&#��C����)�;Cھ�OteJ[���D�C�#�#I�LD~����������w���Sh���ƛ���d]kh��
�׈���F�֫�5:?���&�4���&�E�ѕ���W�]1g�hҢ���}�-�(3�#�kلL��`H�U�ss$��yh6�j��[J�~ֵ	9V�[���f�O�'�O��K���eX��Z.��ҒJn�_ɤ��aF�8C��M��@��4� �n���7��}]�]����$4S;h����Eú��]�5��_JF+�90��r�:r�͚:���s�Ṕ�T���
�l�j��}v2�ݻK����\3 9"4�u�ɝ�\:E~s$Ƨ�}P�>��K]�������2�,�+̻�a�S�ow�rG$O[^q��_0�t�|��k��ނ���'1w�'�row��H:�f{M�U:W�ƅ�"'w�;H�֜���7vp�mR�S%bg�y���J�;�rJ�y�'��6&�]�:�{�ѧi��{D��azU�Z �yb�ۃ�:����'C�[�8~ћv�Unx�Nϣ۠c��_w��s�=/��r
7���gs.����PMfQ��#��)�FP�)�;
�(D��4�HE�A:""-(ꠔP(]�H'�z �$�������]�w_����Y�q��s�>���v���\lUu��n����p�e��^�i�kWJn�b��4-��/z:����{�y���hK���q&�j��|�{G����e@5���mR���ni�q"n?~pb+��cV
4��� ���58�w�����Tg�ON�-@nn�Ȕpt�hB2�>Ι��^�m�c:���f��n�x kr��6��M��{��n.���]��	�^��;����w4������(����?�D��O�?�D��O����Q,w�}��t��������G*�a�j��8��ess3������.S>�.�6��E �M5;ח�fw��<G}����
,�KD�r�䕏(V�M]wi:��Qz˽�w�ƈ[��N�}�<��HS��ȃ$�Ra����
@:e�I.����x���pj��E.����͔p�4(ES,w�5>5S���_��Q��թ.��:�q�d����*�]�O��_���(��.��k��B=�!���|U��5B(��t�X���n9,�U�P�0��f�O���Fn��g�WW%����{��}n����W¹��~��O�
K�����=>����V^<�${�n�۷o��~5�T�P��RI-��um���dP��k��9c�4qM�;y��^H�/^��@��gyp��2��Í�Ύ��ן����.���<��}a��dT�_�)/]�F�r��)D��oom�ඬBH��<QUES ��HҾ���k �=��q����;Z��j�[m�;F�����	e�=��%-�g��V@yG��*�_�П"���'��FH	���\�t�α�[�Ł�2���<K���w���~���'kO�	��Úl�p������Y{T��2tJ���H������\$!g�7v���1�����#�#45��^��@�!�j�5ߏ�Z��A��0z�֤�hȔ`��LW����`���!Ͽ�0O��No0�65���]L��X�ʽ�&?���ի��mi�j�,� ޣ���D�%ni�H�!��r�cD�`4)A�љ�<��n�����3�a7l��(pUY��u�8��"qi9��bBi;m���IF֖�J�?�)�:�G�G�r ��sjϏ.�˯΅���\��2A�i� �咱��&�=����DG���1��_�V�yɸh�;�<D�x��y����It�����0�#��xM,_D�*t)�f�K7op}�%�q���a����m:6|
��1
����
�?z��Z���!G��l�y��,��b+><q���@\}D /}��~4���1:\ӟ�}��h��?rZ)��u��4g�����u)Z_M�zN��; �E~>-qͪ0�>u^X�M�M���Z�l�%&�ż^[��lME�Ѫ��PNvRMJ#�F*[ :#'Kp�?��yq���l��g���$4�1�fu̪��*������N����T�ՠ�'�k���u2�د����[#����jl6��p��+���u�ܕ�A��Q��oȺ���E��L�����?o��JQ�BQ�ZG�
�[�UK�]S��#2���H�����x<�.�8�5d]��{���
�zN
�覻o�����\*0pjE�}�@v��}c R?W��w-�p��v��8pbǥ�};�����������_��y�����/�<k��!��`-���Y�l��dԗT�������{�\�דN׾���6Ɂ����YJ�vk?>HG��sg �0yQn��k�4F$�5Į�b�Gx��U u$H�>�]�k��`�<�c�b/o�D]�^�����7f���������1?(|�:�N2����1��wא��{'جn4��>R�:��#�<f���L*|ϒ5�x@V��Q�k/%4�
�
�uF���'�$��n��A缢zE$T���������f�\C|���P�Θ��#��RY��819���I�<���o��C�XǼAZh��+���Lq��M#,�X�8N� �4p&N}}������-�m��c��+X{A�������>�=�F-����kLh3��X!�����m{�p�{jf���c�����y�BE�f�#E\L�L����+K-Ǝ,< {n�0�Cz;��\y�L����M��2�����:����Ck��}N����������TmJ��h����u�W6���߻܈���1��E{qa��X�z�*35�	 � ��C���}��E�jʜ7�z�LhC"���kGN?�x�&'��+�C��ܷq�/`���
�������y�J�W�@��EB�_�#�&S�����?����
�1F����ӉK����"�&8�S�[uB�b
�T�2C]+�I��ty����,��@�x,@̺��7.5v�/��>* �/%.�>�V�^w�J�#�x)�����S%[|�/��;�o~� ?.�,��&>|�l3��t���Y��������w*�=E���� #��sI�ƽ��FD)9�k�B:���IS�ݻB�]C�W6��;�_����x��r��y+�I�0���ɩ���o���|Ȑ�F�]��
գp,��Yn�u2r�ע�à����K����z��R�,�tEҾ)����{��؍���6�X� �G�G1um%$L��I�j����e�0�X[Kv~�>��w:p�z���ar���p=�L2:��ݶ�풏X�d�q���]�#*\.�#�ݪ�+_+�2�30�r�j�������<G.�~���
oBյ�]+Ei�׶2:�z�!y�P�����k��]���t�A�TI�����\)o�{@\�F~����2��_�k�^%��(v�_�n|�-O���H�Mhs�z��Iv��}q�k ���mÞ�	�]���@�؛����,�w�Q�qKaa��X*�R��<:�J�S�`�W�iK���B	�C9�,��������D��'� h�o�TI!/X���M���5z�ڷ�/�Y�qĕ��\�C^�����������ג��$S�ʹ3ل#V��r�O�ؖ�p�w�f�t��}W��S�\�+�7\�N5���f�]�p�"[T�D��ۏ�_��uvv�f������_�.���{�a���W����>�5�"�KZ~���J��\S����^�zspГtGW�� 7;�#xq��7XM� �i��D�F��u+�{��|����[����{��Pp��J�����Z�?��=���4)���a�hz��GD	?ݺP��	-�VO/d*wM@M����
<fBU����eW�IYɺC�1u��S��������5���H�X2y�5V�@޾�+�. l�5�aeƄ[n5aM4�Ɠo���S�q����|�ˉ
�(Ș�����K�Ԉ��� ���/�	�v�+bkF�Q��#?*�Ԟ��vШ�~��|�����xA��R�~�T�^/oQ�0e�����Ƹ��������\�91��A�No��?�bR?]Į��)&&�%���e�U��ѽ��3�2���$�}1�DQ���[��6Å3!	9�o�6�?x�T��G��e`�Y�-+,999_�\G�͕"��.���܁\ȷ�X���\���Jy������Gp��L_;��y88�䎳 n�����*K[��+/S�_���3n�)�K��H�[���?r���u�#���<V�k��s���2�(����B�Vl4U��dqa�3�
f��ʄ�X�$;�',�����yxr�RdY�54�D�>����ׄ����O4ϑ�m�G��"��ɗ���P��}C�Q��sؔ¹
l����A��'ob�pw�>A�q�7��{�8
�hi���8A���=�d���~���$�Y6̄Y���e�^0g��}�-�˸R�ޑ��m	���8g�4�ח�ó�h�3������>7��>�o�9CS��5T�j繐G�B��\�3ԝ�����`�}M�e#�.�vK���*�]�������u8>F������e]ԿC��u�O�L4�.��H�*�nޠE{�F�uӏ�E2W�
/�+X�	R]��K�)�B���W����u�?����7�ӝqoI<��v{�e+�'�x�VU��{�h����=��:�eQWV��R�bg��vѾ�Uh'�n-\�Q�/m�
���&]f*P����8.(�����d��:3��	!��â�;����7X��>r�~Tu�=gb�Z-�>_�["H�n/�a���K�{<`��,:o�;��ci�V`�,�h*�i�XU�g���^�T�bsr(V�D�����U�_p���K��ÂABe����f�:���q�?�V@��RQ�L`na�ix@�Z��ܞ�����g���.Kp����Eb����]+kd�vz�����,�>�;�I����p,��Ç���]k%��$Q}}}���:�5��9�E�������r���Q�t-{䉵d��x0���>x�<K��3v�����0��m�� �����y��䃔��&뢗�'�����i~F9!�UH	4�Cu�1�� g�濖�L��؁��Xy�r�\a�V�Llnn���t��S�N�-l���'hӷ
�� �;���/����!����_�	N
F�zf�����dt�cFA5���^�UfA�Zu�9)i�lA�d���WTo�	z$ ��F��P���n��|�����B`�N����G�Xg�dLyy"�>�wB��߇��\PX�)z���2kH�E��Ӧ�;��#�:���t}�6����5��Kd�����}��X�L`��.��~��P��&=NPY�N�n�,��/�|���S/��g�/ʮ�vyX���]{b�滆��3T�d=<�$�Xr?��CF����gryX�ԙ��i�����*��0��e��\;"�ps;j�jr}Hr��%�6����x�P@����i��=�]��pK[��[J2�R> 0�7�BKl�/��/
�K_��	��t��C�LNNc�c���q��=Q�󆼞��^0��Oy��Vg������ e�^,N�����d����.+j/h�Nq�6�U�&���Z�fbr���`�>�&��lsFe9�X����[����5)����Q#�|h̢+� z=i���3.Z�<11QǔȨ?�4�� me�p�IS��
S���Y ��".`��ԙ��\��ҏv��_l\\���n<;P�Ԕ-�Mt٠S��(�������շ���`N͆�_������q#F%4?�:UFU������rz�]���~��\�[M�n�g���>`�S[[[��;�����Ph�67w��7�39�-���
���CX�3��yh�R��j��H�tvvf�'��X4�<`Jj����H�?�+F����^;pr�����e�I�+<]+ �	�zzzZh�t�B]���@�%SiQY`ٲN�\��R&'ݔ?h����:]�V� mu٢�f�&sh)�fK{�=<��P��-ҐM���N�@�~s�5����qxju�K��h��lv�2L�Y�ͨC���{�3��
9��S ��(�7���_�+oI%�b**-�X��(ⶵ٩I�#\e��d��u�(]PQQ���KNO�+@00�Ծd��|�UN��DGGG��V��.�����)���n�,Z��e�nL|�tG�e��fuH�����8���>`)\�کEq�F�E?�����Ō��f��i��"_���(5��׆<M�u��b�B3���<�C�j}�x���އM,��:r/YF�\"��"E���=�v����|b����R�=�W�ta�޶�璋7z[��~�y�Zٛ=H�^�C�o��)��s���=3]���_w$�;o2p�8������wށ8����GyR;@���v�ꏷ�99�������/�Uȳ��>������y222+3]=��'`���*�����CCC��&�}��:wy�?���9���������_h��K��P6��&ݴ��ٓ��̃��%c{�K"4�Z���4�~	B&���1rUN�h�td�#�GPs�MH�3�%�Lm�jӛcb ��q�t�����c��;��]�WٵJDPWV�+��.J=Ӆ?Z��N�3; �#��!��1N��iN+�TZ@����B�vu�-7������k����p�?�꯯�N��y���V���o�w����bS:7��Im�����M��D�����a�����_OA?*�<;��>�f�_��'?I�x;9�Ư��S�c�Ϝ�{7E����W\��h�	xv��ġ]��rq)Ĥ�9��t�`3G"E��$�����S�!�>�D	�%�B��|]sՇ�<����K���"���k���p1���� ��vK.v~�D���G�OS�ͪ��瑧��9�iԖ�Vw�,,縕Y���r������!o<_	õ<����+��������n�D��7�_#���NC��V��i��|�n�m��˜�6q�&����P���Ē�.�B9�����΋@7�!T}��ƊCW��Z8�۰�&F��b���\���e/�;���0a�6&$�"]\\ ��(,\H�K2Щ=K4��w%����&�%ʆ�25I.�;��U���#=�VB��°�F�^�ТT�"$�z:�5�:$N�8۝�a.��i�n�C�u��!��5���bJdVݥU%R[���s-���}��\6�	��!�����՟�yR��?_5��r'�"W����=�:İ��򻰨�/[��g��ot3�55R|!����4%u����r�����`sV�>�p'�Oۀ��M�ŵ�!"�8w\1`�<�*������g��W#�^(�k*T������}q�%��w*����*ɸ�[�Vi"J����ݔ�aQ��0Y���ɧ�a�E]��Ο���	I7�:�����ܣ�G�(�[_6Z����X�{j��y˗�g�Z�U��cw�:�1�%VI�G4:�p�
�vy���ĕ
+;��0i�_��Z����6�M�ǒ�
/�<��@;�DݶBM�U_ Z��՚Ҳ]�>�2�amu=!;��1�g����/5'�ͅ��"=�s�k���v*���G�c����9�<��?��O��s�d���m-���}zG�e��02R�R��}�*��_��5q4y5aC���G4��R����e���W̌����������#oF0����~��Y��@�~�P�vrPk�V�q����|
ћCB�~Jh��GO�r��-u�PIԅ��K����ِv�Z<�ʚZ��M��8E��v'^�48�@���JXc�	�<2"d+�c�����ҹ�4�$�{W��z���>}hY��R%��5��~�q�h�Q���k.�y5
��wv�W�g����ɗ�%+]"X����.��MW���R��3vp��t��ދ���T1x5Z�h�n]u>D4�צJ�ۇΎ+*T��\9���}���i����|�|����(^���s#Z�5�]�vэ���ĵT�Q��]���-�JL�/u|q��dKn�bΌ=Ito�j�S/k���E�^Ws�:�)������UEBN<��R��z}�å)�҅��i�7�U��o�opq�q��e��=9�NC���mP��o�󸈫0#׮È�O� �y��+�ֱ�/SF9���c}!ޯMרH�`�բ
9g���(�Ό������K�M�|q��w� Vr��$����8i��ܝ�;��W��!���@#~^���
ǖ_2Y�C�7H��d���uk�B��X��,ת��{�l�K�W)k�mPͧl%��bdi����ң�LPDs/GӪ�t�m���m����XH�v]�&����wS��?7, �=�Y�пw�/��W'°K�J>V��>t���O�	Q	��+��oP��l�Ǘʩ.�f^�(_ݒ��͂۴���9�}	��{�*��1ۧ$�g"���XW����Cj���9*T1a�T�]sv(	g��R�¼h��-\�yA~</GfKO\N�y��O�0����%�cɆ0�A���Z�����G|��4 �Q�W���q�������=y��e�zf�I�\L^jG��\B�Y( /�{�J�w,���	o�'���t��g��j�M��MT���m'g*Qs�6>��"�ǈ�xo��:����sTH�W�l$�{P9w�[�U�Mc6�of�Q�𴮾�Qu������_0c��+�/V�����[�9���l��G��5z*nI4ή���l�<?3��5'��:�n���&�B*��e)�	}�#���Zm��WI^i�a��-�+�o��U.仰�u~�;?ZC���Ĥ��l�
�D��#L`{�s�7Ҫ�b�}(�4^k �l�'[�l��\h��$-Qo2��T6��oe�����+����z�������@X��-�8�]�i�\z��`x�3^#�]Oh�u��Ls�r��X����V�#�w���׈�\]e�H8��QMu�c55dlQ�㫧��)�V�p��2k���X_���xZ�o#n�M�Br%�$�ƭj�V�/���r���N��&�^���mw��*/����M�x�c�cx���������7ڙ���.9������a�k�H�å9/�#p�7&ν�c������h�	o��PO��S!�҇Mn1�B�8W�RH���K>�_�Q�=�׍��Z;#���g%�G��l^)V,����-��yiɳ`N���Bn!G}���15/qCy=&���4�����dM������	�{R�f��Mѫ|���u�t �`���OA�9�wh�P��8.�g��{��h͗���Xʩ~(9��*�u`I�r	YTekd�qA�4Ds����ͬ���	�=�nհ���� 7�{���BU��B�����w|�gA�:��D�l#��t��CIw��ê#����β��Ȋ�e��RM���v�q�gc��c4�3s��^��b���h��n\X�@�5&��F�/�5�����S���ޭ��f������=xr��[���w�i�8��61�����!��6�%'_�kظ9	kT���;���plX8F?Y���9��Ԫ���P���)1{��� ^�YSs�B���2>Y�󎭭�y)-P瑘�m�vcU�c��G�x�����<�q���޺T�5I���Q1N������;����k"q�.#�zzzK"���YQtC7�4ٜsaxm�X��Ƌ�J*��|0Io�F+WԻ���z4_b\�����FH��f��������@1��:��j$Y�.��+�!+���c��ѹ7A��!5,AK_]�\�_1�0!�Zc�q
1X[�#�&�sL�^`Z���)kw�E�W&ʀ�WY��h����,����%����j$�ZV��x�$Er1����.���[#ۄ|�(��p�Y%a��Z��DZ�g,`�q�ڧ��.���^t#�m��'\�4�<�e�
4�<ahZr�
ȝzz�]9�)S,c�(F������H�<�-9hX�aA��#��lT���oe:Z ���9)o��f
X��լ��W9y�^=w!����%�O��G-��8L�����ۡ���-�p_�3HC�� �)5v���9�CV�+ҽ[�������2�S�u�QUz=�x^R�Sc�O�	C��u��~@$�ߕ9���<�?�R�1�	4�d����8x>�Cn�xn��l�xt�7�X�#ӷ���Q�Iŷ�ͨ~mw�ʍ;��ӡe� ����_�8C,���$�4(�V'2�8�hiZ�ϔ��� ����]�Xl���[4j�>��]�hğ�,'Ʒ���3E�+X��ي��uu��k%���T�;*�%��#T6A��NC�߰��kZX��\j���NL0��`r���Ṃ��'�@�d�����\�Z��r�v��%o��s6�g=���K�$,�ñ oБ��cG���[�l�<�#x�y\�(��[��j�YR�b������m�@B֭釋0�z�e�j����ܱ������)�f���c-�<l,Fs$b��7����69)�	�ל�3�7�1�T`��]�.{_h>yQG�2���Y��y��.��쒳��#�|/K�]�cā<����y��
y�~�4i(�@bg7�rYG��N�r�զ�e�<��E^�䜈J�=6��E�o&b���C�[_���l�a+��?+��d���v)�r��k� a9=�Q�
t$"��	y���5�g'�ȘU�ѵ���0.����f�eǎ����o'?C1�.j�o�
T�4켒e�� \����3ɍ��4ߚۯ0�����=�Z~�ϣ�J�0���A�E��Z,�F[�P�AU�؁��*;�P[�Tp�����٭C���)��������Kx�\�ĭ��܋\L��9��ҷ��{�Q\�ّ8��;�Y��<��T+�a�ǛҷP����I5`��������A���v��کk/��o_��Ӹ݃�|T�(ˋ�.�'���ߏO�\#�����{���/!�`��{�a=I���KA��r5]"��.�FJƥ����B~���U��Zv�Z»�\�8w ���U���9<h���c��ނ�ԓlmF����	Une�������W�@!�kڂ_h ي�ra���03/��w�����{��U� D��rg9�D�~2x%��������@<��T.�g�%�/L����4�`��S_-��^.T���ު �9b�8��� �����tՙ�z|�A��*r�4u�7g�Z�36�7Ns�]f/KK�X����2i�o �xy�d��0[���Q�����L$Y�JG+i��EP��9t=���r�k,޻�2'�9݋9�W]ϧ�`��F�e�/�:a��z�a��Y��w��5#��6���O��X|6��=���θ
�@��Rt�W6р ��Pէ���٘-f�����bV��Ǐ��ܤ��
�ζȖh��I%��#����*�PY��6����X$%�{��,����R��C��`zV�G�b�:�1X}۞�~5�4)XSs�]~� �|��k6D��,��R�Hҡ΄Zua�@�D��amHUE�9��?��A:�*�hQF����^�a�����@X��_f�z7a�k����ـ����d��D �#�h+��0;+y�tLP��֜��������0���.�w����m�m��}@�>���ʒ�wu�Z1����.�[�W(�l<���?39��R�j�{���Jl�����m��׉�%BCbZ�AM����D��bS�*�u�z�V�q�5MBoRԕ�,{i}ix���İ���~��'┋Ͼ��<���k }�j�Y��WGA7�݋mN��?�M�B���[Z5!�4��^���9���`ԣt3������0�z���a@��P\��bsG�����ʂ�k��H��<٢����`xu���|�Q�R�՞Ae<=3R�&�l�G���}Z�j�M	��d�@�"��Ճ�CE��#��4ݮYH�K�T��zh�[�J����(�p���7R����*��m� ��17M�Z�H�2am�O�����1bq�$mc:G�Ve�sd��."L�G$UWc�5��4��!lY�Ӆx|)� )-�<|��ǝ3"Q���C��[��Lu�B7�6��a5��Nꌊ��J���a�4�3�uQ��bQ�yM�e�����f�95u+�x�����h[Ȝ��㒪��5ԵӶ[�Z'������L� 4)j�w��T�J`������1�2£��uO��Uq�-T���Пcgq�;LR^FA]P�ܝ�Ea���[7��_L̟\hԲ?_m��c��EGPO��)�h/�*?�GF=��6 �ҡ��ߪg�y''?��]6��ز��73���*"�����1+_O�(���^�i逭���/�h-)7�(+�����+;PR�.���Ц�����7m�^~���q�7y�j��X��G��!����?��M��vJ�4���wu4��C�j��2� ��>t��7Q^@Yʻ�ӡi|��v;��>J��u�OQ3��5sV�Z [��j���P(����
br��ۮ_`��vKX�C.�Dc�gC@r$�IK���܊��D i�ޏl��>�@u��"i�/`�k�qg�d2��n�G�j�5�(vv����C,P����Q�@�5��	F�7�k��Ҩ�v�A�?X�vg���/�U� -_Mwܑ�7��op�����@��u��	M�.���<�ܫ���5�)���F�NL	 	�(�F˂�2�q�G�W�4����0F'48���H�`5��V��YTl��[���Tax!Ǥ�)�����R��(���?RQ`�>�q�`�a纼��]��.�՚�p

��J����l�����+��/\�Ҿ����L��Wy��H��Z�R�������J��ƨ������v�+�[8U�V�Q��)/!=�5ש��N��;ŧ���zm.�L�oB�Ӊ+�f�����A�l�,��3�i��ã#��WR�>I�3 ���9�$�h͈��O��j��VZhC����^~U���U����ZH�R�3曄'V:�iW��}&�Y��Y�^,�,��ʓw��
l�L����G,�l�	�1bN��&X���kX.�?$x�@b�%P%]�TO1�����P�ˢM�k!���[�^|�;<�I�h�>p��͛�;�U�RKv6�ޗMO��yj���%�K�.cP��k���
���X��]u@P%���c��`�P�%^ JH_�N/�f%�i�q��Q��,O�q������+Xь7�/}��3A���iɕGF�}F����S��u��rer�$y05E���kt�'MF0���l�F�N�v�p5�l���.0��:֬�S�霐�ˍbz[��bH�E|�^	�c]�,P�3����6:��R�ԟ&=��ZF�5UC<�֯_��6�Ar>}u�-��1Jڇ|�㿖�k�Ԣ��ÏT[}��&����4�&��yR�;}ݨ��*�Z[�e�!<i�+P�P��^*Zhw�.����[�f�M�識�1A��r���O���T�r8Y}�ՏP
k`�@.��q��z�U��(f�'�/y��<�_���N E @i����J�אռ����K��H0�m��x�����5#t6�L�
V�淐����8Uc
�8/�	X�.1��h�%4�Eh���v=����g��2�6�Թ�q��=L��j�FOC��4��N�Gծ@I@�@`@]ZI�@g�ݾ�.�R�F!շ��V�=!�#@�^tC�����ٍM:����By��$�O��(4h�n�"F�M��N�M���lm�[E��z�:��%��}Y/��ش���9���R�H���gh�!�t�w��8�D�fc�w�q�hrv}���8�Tt�q��>��V�S�>S+�k�	�Mvx�7֥`�Ɉቘ������Q��U(�!�I6[��]��c5��_�ʷj��j��+-�ǫ��9�.>�幒��s�0�YB�JU/�K<�ڄ^{{����(���Z���4����P�M��\�`6�OU�R#�.�+����©�c�%WS����,K	�m�C���L��U+*	4�O�Z?�|�8��_w�
��+��\aD�I	A��������ܒ��|u�E~?-�Z�Bu�6�A\������H �/#s �W�ďjjO�x�vO��k��7���4�	���C��ayD�6���Y�d�����'Y9���q'p��z��B�i~���S�g�33�x�T��%���{'�!j� �O
��9�4�l�B���Q��V�w0�`���Y��eM��٨g����Қ�Q��'������^g����Åѣj��K�=��j�#HS�����"�!�+�;�N�`W�U���Ĉ��D'���-�r	@�ԓD��gG�B�\yWԳ�t\����s��~cE���'*3!ސ��4�pѤG1�8u�^���P���!��e�e�k�a�9���þ��l�~.Б��zFZ��T]i��+��τ�|�
�R�I2alY�_�'��?$1 dI�92n|VVǨ��-W�L�p�TT�)<��xT���]�bƆ.�B�JHN)We���{�%򬩥�i>^П�E�a_�Ɖ,�Bi`%��ƨ��U^}S���oT_�{��7�J���-Z3��{}�CYAt~!|��Ja��`y�`�R`�S��]3s�$�(��֯_>�6
!Tױ5aa��1�4ػ'g� �t�_̛�=�����v�u����v����gl@����1��*����ꗆ�M��0�[-�lxA;\���`ݼ����1�|p:H�]5��y���yŚ`��GkLô�a���O��m�k����13JқC�Z0G��RG��e��������D%Y� �77���gxAmWk�!���/����g�s�b��8W�|FY��7�%b���
����X%u��>,�֍�_&:�7R$��zt񵒊
g|�u�=䒾/=G���������Wm	��=�ԾR���RB/%;�d$�r��s��JO,���澄��ڥ������;F�`v�������/t�j��+�a����{���_\������_�����g������V�Ż�7PK   �	DXd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   �	DX�Ƚ׌  �  /   images/9185dcb2-65ea-4de0-8d42-42cedb1b5634.png�x��PNG

   IHDR   d   -   X���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��\�o��ݙ�����uڗ��!Q�Bp�D"��h(U�$B�F_���?�C�JM�!-�А�J�(�U(I��E�|�^$k�w��u{�ݝ���?���gM|}?~3���眹3'֎_�A`$�M!p�8	Q����~��Ql18���gv`��ű�K�Vr���x�p�z�3���rW�y�4�0Ɲ��t��=�r�Ҙ�xq�!4q]&��:׸:/s����Թn�?V̕%�p���:�+3xg�X�@?��Ⱥ�qO�W�t�G�����X�ѳo���Ij��;m�I�Ae�ŰĠaä���	.���'�eV�	C	��h�*��2�z�=.�q�k��I�%WZ�A�KD����rB����'H)��8�{?J����>�9���v�4�'���~��.��7�'`��9F+ o	�'�!p��/e��!i{?�CP����Ij�Ҹ<즺aj;C}��Ǘsݥ��N\₱�ߧ�$ސK�\��G��	y��s���׸��s��%\�I��,� ^�cg���CT���;s���/��e����2f�f�}x;����Q���r�����2	��b�\͘�#���-��pb�w��u6�S��;92���&�}�5L|�,�a��ʚ�K��D1p�eM�H��ugDq�ߣ�[5.W�z�D
!����	q��MB\s%��Zs9ߦ{�/�$��b	ӓ9����M%wk|ao��3�=�)㭱�I��4Me����K�_�%?�q�<��5'��-����Ү_���W��:�of?�˸S@�w�ۻ��~Ϋ�1\��K�
�^=e4��"������W]�r�\�ո�k��書��հÛ�����$����ǰS6�}�������>��ذ�)���Ty�"��])����ZMtXT^��s�V>�q�<C%C�u�2�~󘫕���M5�;s���R^����D����}�s_!�.I��VH����k!�){a���2��0ڔ[���̵��`@��XxL�zp�f�S�7B��"s���q�<σ���ҿ�P��J��h��Ȝ���g.����U�^}Qx��t:��C�Z%�d)�jдЛ�s�1�J!�H F����R�����Ӓ뺈q��U!�M�#���c��"(�Bt��]R*��V }�����H'��t��Q!���xUH~&a�����!١;غ5 CG�4�O4䏱z��אi4)D�Ζ)�L�8:$�U�vQ������:�Gx��x�.��~���n#���q�EA/W�W�H��s��������/�]]T<���}t��.��j�G�E��WX�_�|BE�
���Y�0��/-S���F�]̓����@�1����n���~k��j�ل�C�ޠهđ��CW�c�+��+���\�B��T����8���u<6:.��aYC[q��Z]C�r��X	�z�Z�Z!�Fcr=�/��Ut���q�@�\Ѱ���\�d�\���r�r>jp������!�=w��B��B����`t{c��	��겻�GA��lZ��v}�m��_�Z��v�qb����/�^�B(JKO���'a��iw4���������~zHي+ڮ���E�S>��W󉞻�S*;e�d��vr�-�+�hVXG���f䫊u�S�#�J��Uj�pc��mw|}���l� i�!�x_~=����oܺ*�5��S������q�8N��\����MW;t}c844��'G5���!����}yB����a9F{(?"�_�$9�c�3TC!���
)|�B�O����ؗ��0�W&�RxT�R����s%v�iѥ)��	^�U��=+���0-zJ(���/����R	o|�6��}� �3n�����=zw�G�X�ξ���z0;���<w����4^y� Ο��R�¬����i�C�8��y,U�0��UI�c��W�1��u�Q��\�����p�{`�OO�0Br��V�u�0���\�=�r�9=�Va2^��ͅ	!�sZ4+���w�n������ة�jep��!b�~?�7�՟�{PiѤ ��?�(�*��    IEND�B`�PK   �DX*�e#o� Į /   images/957f05b2-baab-48fc-bd29-824c654b1c09.png�eT�A�(ڸ;�-8��Ƃ'�����%ww	ww���Cp�Hf�93��u߯���1_w���j�����%LIA
�  �IW �R jD���Or�7$�Z�  
ΟH� x��hJ�HK� �v^�C� �^������0  �?�?���0���
�NB^����F�O8ᵱCA�^���
��K^�y(�_�v�?.Ŀ�p������������ dr���8)���ٸ��9^��r�G�?�[9ҫlh.檚N��r�ƶ�,�`[#����_Aa7;CcK�����Dy��IIaQjpɳ�۽����p��x(�{X�)�����_	XC�)ܬ�l��@�����Y))��8Y�(5_�~o� ��d�dac�p3wR
!S:�M���%�I��4sr��geuuueq�`�u0ee���ce��̯̎�6N�n�6�TH���8��������ֆ�O�����	DI�:O�_�Y����7y�Z���n�v��,l��֬����I�����Q��ªq�uv0�H�@l���������9;X�Ul�
��X��:��`�7��o&05�����U��t271�_��g�p�/�����E�k#~q[c�?�I��(���������@ ��	�	3;'3����'/�	7��k�c���R�6�N�6Ɛ?�^GX�_���� |<̼Ɔ&̜l�t����y��l�&\\&�<�BB���5*��U�?�����^Ip�9y�yظؘ9�x��!`.fૄ�l�`NC�_R`c~I[k�Ww�[�BX�lL�N�18���4����?#JV�N&�^s��l���?S���'�?�d�a�ac�bg�f��}}��:���5�P���g�8�:�J:��e�/=��;@�lTmm�@�����=-��P`C'CqC'�+���|���|�?���ۂ�M��������?������ߡ�
���t���ѡ������P������)c3CS�k�`��q��E0��p�p�q0q�zhb��g���`c#n��h�w*��&N��Q�W;���5*�ڊ����b�w|W3��?���d�#pS��SY��V���c� �K��S�X�Y�^+!��������&�a�&�a�&�a�&�W1A�����u��zT��y� ��H����e�#吨%
�X�4Q`�8��wC2>�D=�a�1�3����~$����å�i�jBےܣca�A � ��PJ�Q�V��v:�������.ˮy����~�4W�z���q�󮴬f� ��U&Q�[�:u�]�ｏ��H�R���s��$���Ri%Gc��Y���S(�!!���2�N����660������H���-Ro�.�[ZZ��KcO�,��vt0�]�Ϙ퍦�ͩ�L͖��U?�u�����Mˎ�
���9���M>�y[�P��m�z-iźd)���2_�O)�	�4���g����Cy&W��v\FKӇ���(T���#=H����	(���e}�,�ל'@����J���6�N��"E�[��Ҫ��ЮN\�!]���H`����È`þ�;���Qsc,�v�FQ=� ���kH�r`����ͺ�ӳ_�"���t0xv�/x2�V��9&�Z$�*��s��8Y�
�3�q���ii���J�*���|�
+s`�@���_=��h���j=]�1P���`ǜI��7��ݍi�w��}ϥ�"�;�Cۇ��J_ȩ���_�jj�����hyw� ����K�G-���e�I�J�I+�%ޗ)���ASrM�� �ބ�7=�g9��o�L�5�OC@�~��Y���q��+��]�}��>��Ĳm'h,E(�e�Y��%���]����e�G�`k�J�`�p�_�UU@F��?ux�qUdy]H��A�TN�_gpE�8|^���M��� �R��<M2���sݖn,w�\�v�~Px!Y� ���'�KU7r@���: `bHp�MY;��2���4a�<ƭӿlq�Ѡf��k��|��������kk��]�����'hޱ�s�Z�n����#�t'<5�%�zd�;b��>�[����"�_��TS������ҫE��oj�Ί��a+�����M�17b��üZ鰉)��R����Q�M�p	`|L�h�b�m�^.8&�̋<~;x�ɻ�+@��E�1�.�{)x���ّ%�	kϥ���0��c:���h����౻g�g���pVd���;(1����55- �z�g"��ϱd?�����ں��^����f&o�rhs6l�����m�᭣�&l��|,��9M�����	�����ʕC�� A���QB�G�c��wd�:3,�����/^�&0B�C���ϗW[��)�'��Q.�޷
��4��g���ު��A�{g��B��[+t���4����+;��3X�)���}�{c<<<xG��A��nH�]4��2�;y�d�/�&]�}�06bq"(�!�v>R�l�.,���-�ף4�~9�� ��b,&�߹n�U��W��>�7����~&��د�|��]�2'��q�i�aK��*3�l*j�Ub��9����/L�!����m���M2�l�uGi��b4
`����)ǊF�6w}gE��g�๎�!�OG���VM����d`��ş�E��wE����y��ֹaߴ���gM��{t��b�� F�y&�ˢ?��)������K���tz��y���2�T�uٚ'����@�6G�]�|�Y]}I�Od3�۶a����V�zZ�M�D�#�3L�8m�Ob֑��r�����mB	ܺ:�Y��P����^k_b���kz���Uuh�=�W��(aJ����Lc&��g���� &����K�̉f��T����'qGy��
�BU�sip�Ҙѣ��E�CL�J��!�߅��y���/�t��h�
�5FxO�|rY
�Y2%Z�~7Oy��hi�M�[YM�k�k-a�Wi��%oߺ��Ky,|r�r`��t�~����Hu�&�=[t���v3��z�-f���j�l^? �!�;�/��Ɂ�v P"�[���c@G1��>��=�	�(��t],�PiY�
�c�bQ7��VG7���%U]F�����G�t�P�h�M�I���W8��\=�9����v��ݖ	�]���AS=-�`�;�}����w1%eV'��_�5��i�/�w�9��{��.:dm��gB"�8�{  �M��=���{i��7Z~��I�!�{�H��>d�T���p����F�FϦI@[��$~���=	��Bc�$�WO��N�� %�-�ԕZ�S��m���A��ʝ�/�k�5�6���mї!l���O�-g=(���/m�����]�y�2�47�����X���/q����O�Y}D�}Ǳ	RBp�ʶ��o
�P���~�8��!AZm�g�O.N�����k=����u'����aat���FJ��=k��g��8)���xh��+�Z��.f�)��s��h��=�������-DbB�E�Ev�d���>�P*�kߘ�:[�^��ϔ��"�ɭ���aYy�U���d���'+2t�5�5�����b����ܚ4-�/ZL)�w�R5�@x�Y��R!�%�w4.�7ޣ#}����S�Q�ͭ�.vv�҂.r`�K�x?�v ���s��~�#�e�a�Vg��H����D[�E�
����oc��x�(.Ǌ����S��h�LF;��l:��MJ�0|��ܞ<�Ka��0x��8�a���>c�z٣�	>�P$�ټcԲ�"Q7�~���3�6t���'\�a��C��9���ۇE-��*� 2F� ���kM�G s�sd������
R��?�0� �Qx۰��Ż���:]������$��{�"@E�tt�;{�T��(�P��4Ǵ|�Cֿ<�T����c�wRgj�/�`�;N4�&�vUV׏_nz~<]
BsߵH<K��;��J^0�K��L�w��#��f�Bq�k�X����?͈�*��{�z\/LA�.���x���dw��A����u�Y���R�=�F��uٽaݷC�v�YP�1��ܾ*O��z#�˂��-�\������$��� �����y|��y����\�����2q�� �U&y�P!��%��9���1��k��E~��Hߘ6�v��lM}N� 9adD��u�o� �.��R�L(e�����<�:��t���{pl�)Yl��b�i`k9b{{�Ԧ�?j�<T��)y�02�vߦ�u��9B�.����Ǘ��[�� T�ǳރ���=X!��"2�Q�&7z�
���,�#<A�b	�="�cD��$4�X7��LS?p����^'��h|##&A�"� n	!�VW��C��S]܍|ݵs�	�ǖ���%x�ߍ�͗IӸ��l�NP�����wQ��R��� �c�D�Ez���;�`�uU·�/�������A������˭/��L�	8`|��(;'��<RW2˧��4�
��3����ʻ�{�\$�	��ß�Z�C�c̻nk]��g�c�	P3��7�pv�P�^�*�0��C���S6H7�uxV$6��=�.�=|(���H-�R0�)1\�9�*��4:ގ5=��EF��7{|�oɛA�3�J���ry�7M�T���@��`@[	�W��qJC��hw��	HHҨg2�?�"-�t�:����o~��̏�-7͉&�����B����'�V�Nkח���\�t��Kg�z�J��nMl�����봬�6�,j�3 �$�G��Kr���-�R1�Igϛ/c������$�Vv�p�5(Myv����>yK��h7�����FgSB�O�9c�U{��&#U8r�B#��һ�s����0}
t��"T�>����}ؿ~���o'�SG�"L�<���o%'��!]l�JU��������j��Z�nZ%R^(�f2��cw��M�
^L�lv��S#E
�"�w�fm^�޷��?C?h�1���N[�/���r�q�L_�[`���/t7�
/>�tr����ka�X�����|���/���H����Ǻ�Uu�S�?����/Q�q��59PN�~�y�3���e�qG�m��mAn͇<�f c7��+*K.n�$�Fs�{�\���Rƣ�V�M��0���K�J�Hs߰s������1*�2
Mv��p.�ε�!�����"S��R�L�U;H?�+�N��h�@��^��]k��7���/>����l�zL����'�d<V��f��AX4�d@�,�,�D��֥2A1�����հ��')a���o&C�0�ƪ�
y"���~�n�u�h%#��cϙ�7>��кRk��z�b?��|R��ދe��#��OA��^�N@C�DV=��m��¢$����|�~�����R��`@�-���vrOT�v�/-�GOc _��˙�ϕ)��UEr����5~߷������h	�����G��dGɰ��o�W�����mZ�:n�+��)D���y_�)���7k�J����c����n�;����0M�ƏWq�ݧm#.�LJ��9n����IW�$%{����!�C��jt��\E$�W��%�?v�x*��]ɇv��Hƍ.���+BJ���|e���$�����s���"�)�j~LX��� 7�~��		��)�_�?V�\�3c]�}�P�ҘJ��hN�q��aG ���g)����}ƍ#1��Y|u:A�G@9��������]T��Mu4�,*��}��
�W3�	��v�	�3Yl�Ba�ݩ#��W��Ńm`�בa�P�ʂ� ��c[���-(�zl(��Xfۓ������=��o��(�~��G=u��u�`~���G���	���:��O*
2#�GuxǸ��.���j�2��FB�E��z������*�NJKJaJ�@�f�i���`Β���v��"�]F��L�q���t�j:��h�o��p@�� �;�pT�q�(-�A�}3(G�A&{?�ܑ�M���)���б�*�����z<�o��t�Y�t��J��ٍ����mk�/H����̳�k���s�[V8�� 9Qx?a��G��B*({��b��\�a^��s����rb=>W(u��~ f)��������)ō7��`
J�ыyH��+���Ck6_�EU��R�"�Ԛ�����n		���vd���*�þ�ڐ��F��i=������?����uB��^f��O�<2o�C�f��q�D��3�,�`:S��F�/��E��v�vd�?¥��˄��\��KAu��߮�z+����>.�s� ���a����ط�^S;y�7��U�fҀӳ���9�C�)G��h0����?ɒ��*�Ub�z��y�gPڐ}��Ɔr�������k�t,�嵔?� R��
R��N��Fܵ��\� �>2a�2IO?󺣳V�����U�p�_���lNa��< !��}:��S
��2	x}�ߞIyv�
�C���_yZ_*#zs�օ���f#�9Rr-���̼î��W)f.�#�ev��` �n9eagɟ,�B��o����I�V9l����	;U@��Ħǻ*�`���P#d~(���ɾ#*�G��A⮿���/s�<����'�՚����ө\Bڔ�u�̂Bf��ll��xe�l���ݑ�_n�:�7��3��So��y���)�s�AD���}�n<��ѿg��~~+����8�t��(U����o6@�:���6I��,)���9����~d��{c�b�C��/W�*��+(=F��B�h:�W"�g^��ʏ�:s/��y�~��6� R���1����K�:K�����^9׼�t�fI�-ڴ�0��̱����qd誁DF��j��Rkf	O0
��!Zjs1���^&�C "�`^ң�BO�����a\X���8�	b��w����&L�@��R�ލ8�!z�D@�� �?Z��3T�f���=xc@p{�l�dc�53��O��<~���y:-ͽg��h��-1!Yz����H�����s�@6y���r�P����ijz�P�k>�t|ߞ�.)k���0x=<d��`q��%3��;��'���L�[sr"�"ٍ(8aB�ۣ'I{�p�<\(קֱ�f� ��%�r[P!f�R*�NZz7������!B&���4�)η6�@�5�#د����u��_E�(�(�w�_֦�YEj��ضs�����$����9MI࣑:M��D p�!sYc���uoܢ޿�=���ɥ�\�y����=��͎6��X�D�]��%+|�4*��D mC��"mΰi�yh��%Q��TL�ֹ�h��W��T�9��>v�G���l��Vl��|`ue����(S�n#�����\`# ��j���F��\ry�6~OJ*wm��/�/˧� �J%�_����F8��.++ބ��׹zˏ]H��C���>?�3�[�}������lf��aA4FS�Sl���/ӂLmKB� ���9��YF�{�#�?�{�P��m��Z���0A{�Ew�׳*�f�pD�d�G�j?���o��$R�oe���t��.-0g���f=!��d����U=$���
�G�8�*���0��C慖����6�����������!���ЎS0lv6�I$v�M�4�s��δ�r�gŏ���6Z���rW��N����֏��̣?��S���������Kv��L-�U����$s�(�/Vq%�Qh00{;��g�4���#���������ٍ��C��C�A�!���]���������M��N_��,k;��=G�t���|���˃c��=��7��R��,b?�����(�������SK��c�P������Jj�}���`is�&����	�q'T2�.�h�BlA���*�g��ְ�B��]���e˔&�6�LƤ%��؝�G]�>�QW&3џ|TN�J�F�6��`Y��d)��2����B�o^�:��5�Kɉ8��$�BIw�+\�������_�8�����S���o�:lzb<��S̤q�޵�W8Ly��MTĚ��e�&�&Bà3�Z�И�dc����>����."L��&:<8.��&;t���.�_�f?��~Ơ��`�-�97~3Q�e�4,�m��ґװ��q��x>`���\ns�?,��I8�}�4��m�ݫ�fX�������%CC��[������=���V�=Y�*���Z��Ko
Yd�
~/o�� Ó��C�ޘ�{��#)z)L@�
�ia_�Z�
�yIS��ǝ�X>��0dd$�×S<De���;+�̴R
��Оe*#f�~��n�M�[ꁕM��l�ٗM&����C��<dɢ�T�,����P�Hq���Ed��i�>��$=:#����;����]|���U�q�;��V�JE���/�����֍S	*f�\w�J��1�ޏ����u�9�f5/���	]��F	_�kƀ�zF�z!�&�}D�b�,}�qTJ^w�N�Y*��nIGnFa���I�%�KE���
��h?y1���c-���t]���M�Ҥ�a�m��2D�ϵ��t�Ï~p�>��V���U�V���lýw�B�f'jO�n����)����2�=����`�\����P�⫖��$��,�5 ��I��#�f���Q�U�O�Iǡ�61�����J�_)�U���ؠ=�3�������l���պ	�0
�*�*�a�2��iU=�EZhof��8�,[ a�*<i�}ɮ;���c�I�i�F���a�5L�J��`<�D�j�����oo�J %�F�T3E� /���x�@5�y�6_M��YkW�5��5IF7���g,��hHQ/�`<;*��ܗ���gp1�l�~Z>����#�x��s1Y�C�����N�l���W,C)�؁?7ʍ69K�A,F�_��#��q�+#*sO����_��6r��Ɖ���ˋ��t��pO���b�i��[L�Y��O����M!n��� ;cE����dp`N-�%�jdp�M��n���ݸ+�/g�N�x7��.ً;+�9�z,��ãe6�����K���9�[z�Q��#Sx;��m:����i�i��;'\[HuX�t�U+Pl_�M��6	 7���&���mGZ�\���ʣ)���EN��=���ܘ3'���>���T}�PN��L*K��#���r:. 1�r�Hϛ�8S0�e�L&Yzp^�Đ+J4��L@q�즳
Yu����e�Ќam>
8���h���#Qcv@9��-��#>G�t�s8����I�;��!�+�N*�sw��r.�>�!.�m��r�T�����B��]��`V�ɸ��C�)i�&%��$������xy��D�o�������d�9�>���Ӕ���"�i�}�����Z���%<0�����Yq+����Ĉj'�"v>(�P4~����oT�*(��Il6hc���u�O�� �>��[IU�j���Q�e7�]�+�l�#��hYP�CA�����S��Ld�~i�ʙmm<��-�8$�>6�Ca�A���/��;����p���v�޳ꄹ��,��ܟJ_���*����LfkpyCΝ%���N��7d�]�BGW���rN;�qbF�1�f�^k�䜿��C�%���k��c�T�ޓF}丗L}��lacU��Zu�q�c�����x�5�	6p,���a����c2���M��0Qj�3�Û���Ĥ��'��&8J�k��ɽ�Z�$��㝭�@��Z��P���ҵ��DG9�/Q�+Q��8=7���_>V�m��<F�4S, ��;����an)�i?!!��+�)�6E����%D����n��ce�mǭ�Ub/���d���.Q���Qg)�ޖ"s/�;��MOݮ8�j�i�D�yvG��5��"B��f��B`2�bs-�	��#[M7��.���'-� �1�$) c����ș!7*��J�<�˘��4�P��7���V��.^��v��F���j͓]��GBj^�*jh�����N�Xy�y��LKK�n�Y�m�^�H6���sY��H��Hٶ#r<J�b�b�g3����U	k�N���`�����t�+����_P'����W���YG��M+��t����r$܆��N��^�T/����"[yA;�L�%Wk�/|OG�_5�+��*~n���\��n9��Vd����<+ջ���ǋ�+����C>jn�{������uV��t��+�*�Њ�چ׸L�b�m-{�iϬ3���r1�X��jM.ޑ�1���0�m�T��~��� �V��q��Kw��t	!Z��R�S!��qWW��D�!�dS!s��8���4�o�!�c�*5P�$0���/J�*(Gi�4���#�%Ǿ�i�N�˩q�ȼ�ֆ�k��K�ڕ�!F�{Ӥ`njp���B�ƶ
X]�5�Z1&���sմU;�mIx�F�*�ܷ�-�'�}�C���h�8�����Sz��*c�7�e�j�{q�;�u	^�����~YejMݸ����x��q�o�bY���O��+~��g�^\HC���g�,ɐ��fF	�',��j��,�;i���+���GU77��1W�,OkC���������grz�k��v���`6�?Xư�j����a��IJ� ��F����ė�ϰ�#4����Αs�� ����V�u/#o�<&�.���d1���A�R	�tM�o1���B�'v�-�����PO�thَ���E�G�_�l�Q3��C�����{���.�[��eB'[���̯ǟ�װ��6��6s�`1[x���DaSެ�����6Xi�*wv�}1*"q�܅���0~n͸#��3�IV0����,�C��f;�W�&�į��L��B_Uɂ�"p~���Im%:���.R*���z��WkZ(��~~������\C�m������^D�x�`�_:�g�Xd�Cx�W���Y����t��|K��I��Y�uK�\6��V�;�+���� O����U�9����]b�N��̓�4�Ѓ���,�����-;2�s�t�tj�^7�?R=c�j��/g�'�'��uEZ��1�F�Y��t���Dw��:Ûô�P�=��j��	���Eڗ�4'G�����\O,��V���|�x��CR�_��}-<��ż���>�������3�l}h��J�bQ�4�p�c�W���ٲw����U}mp�lf7sH�It&L8��3�R�M8���	�v8���f�:2;ݴ� �a�|�済�	�'E���������!3u�'G���w�>;�B�����M���MXĺ����ׇ�ln��$��=�)e��F�}!�h�rqA[ 3���S�3��������T.uz`$ �r'^�`�*:n����6̸�7cv��֓kfI�5ގ#Xy����}~���DC�˴j�F�߹��'� p�ud�ϴ�rPjM�0��"���h��͜�d)��%���i�'ޒ���Zbk�6$�Q)��`�l�Fٌ�;�����q	�T�,U�8����a���v�,��t�V���~]��{�(%��R,ِ��V%����h�K�?��J#�E6g� �6yJJ����~����+g����Z�VN��~������s��Hx_m5~�����/���ƽ�x�"���Й��㶇үӽ�����\�yI�:n�Ǯ����^*���K��iL�+��-��	R�l����Ӣ?%�Լ��*��`�65�$F�d���#�v93'u�QPeE�����E���Κ���oKYҖ���+���Q�:7Í�opG�|��š�r6����O>oJ�SؑTrQD-t�%�F�˒ޥt6c����.�N�� ?��k^�0 0�l�n6;[�O���s�,Vya��1mkw�P�`��I�!w����=��2W��٘�'��T|��h4>:+���0k.�ᐎG��	�G�/�OW׬mv�����B�2��,��j�-��(���槛��h�8��#`�����^�DbӢ!�2e(�Dro��w�h�;�;S��J�5������=5��*�����O���x�c�u�4��1�� �RmL]^Y&`�g�0�r!U��ڈ{Q�۞	O>�뫾�yR��
Z��Պ�[�g�5�т>����Nu[�M����#T���)�B��X��0�R�YGu�3p���ӴԸ�"���mav��*�(<ZJ������
�& /��M�H<T����`G�ڍ�Hr^�+b+eg���U�o�Iǥ��N;+��1��[��������-��1����I4��0���1nh�2�k5B%=t�32�7@^�^�R�$�"�}�RH�6��Q5/�Ǣ��[�6�����I��Kk�w)d~�Gl-���zEC��E@�����dФJm��IM�$�-Ί��9�#f�.�ar�f��ф��,�	�y�d��ˡ�f߆��@��T��ȩڔ�
9v^W�1S��v�lm���y��s�~�5Udr�Z;c��A�&��17p��CÉ��GD�R:ߦcv��S�����D�Gt�?gf~�&I�V������0Ɖ���L��E����ݦֲ����|>�։=Z�/�4<�5ꍦ�JkUY�~���I�US��i���oMP枚V[�DhI{O�/C����[9�+{t��Vef���ծ�ka�j-z:���u��(y0B�����EB�'������u��Է1>EB���ޖ�cSyVO������M噱>�q#�h X�< �n`�h.Y���z먧�;��TN�y�=��%��OO��*�^��z���@�Z�n`���!��ԫ.���3��[y�2}g&�@I
�/��W�M���!}`�����H�l�3W�wӥp<�gf
�<���?�xѢ�a�haR�DΖ�V>4�5��g<6��/��r��8�i�� �ـ��������W3���]V�ӼPZT�H��F��N�e�Zu���ETITU��Ù���B"ҽ��0ܨ�OIwZ���%%^�	��C�3����f��7��9ҿ.Z�4����N}^<:e�R#�X�j�ʠSkR	G�Y	�}�M����;W]���&*|I����4Ĥ�;��Y��u�4�qSd�7l���\�Е��M�\d ��Ӗ�!�����&�'�n'h��8. ��Z��(>e�	�x^�y�	���)	�" �˯�1E��=�_ I�U��/�Z��򥴤ڡG���J�H?��|Y�.���SC��LB�,؀�(d6׺�8�g��In��ӡ�/__�'/)��ik��Q�ݎhA`��1��M3���Lv�>k��ZX{���,���{��^�hid�1��@Q�ej�����ߗ]2lpu,HJh�aE)�*�FGU-G5�1�Db�����j��#�&� _$�r�1h��kg�V9d<|�b5��=�:0���vдvR,��0+�K�9��D,Y����,��垏��n񑹺ݠ	��!�凧��ch�e
4>��HùD�tD����jȂp�$c�\ B��R�q|��w
|(�J�9��e'��n�$�x#� g����ax��ӕ=��Fq���\��}���oX�_nfZ~��~�R��,�0��,�2�@y|��-tU:š�o=��_lB��36��Y}q�A�,n����xs�"{���	H���Ӥ+���+��h]ecqn��<�g����)��n��s)!?�\����V,x=�h�����qP]��~�/܇@�h�BS�9.�»�Wc^
�:�Q6��-�-���i%�h�%�༗)��;m�˷�ǐ�>�t�1hw0NHژP���q3�WG++�V���!������������� ����w�[!R�0�(�7���P)��X
g�#,^砗N��yA7ǣF�ѵ@��A���@{V]��\��=!�;L�Aӝp<������Y�TJ�+-�q[�V�����2��J݅��c����|��9E�J��UX��A* �Z��W�����@Nq�8sJ�/q�]��L'�*b&�N�$9i�`�ܑ�?��q��i�S��l\�f��̚���L�i�������O�G?W<��#:;h���V�~�����2G�	�%������>k zq�Y�;ˇEj�߽��U:�i�ź~��!�a��t�A�nl��dݘm!���,��*ô|۪��\��p؉��\�D�c:��8y�R�T��_:���o~�!%Ѵ�^��,y�k$OlrV����z�M�-�'s��5Z�Qpt���y��)p8٘f8P�w�ӭm�A7�6M�Y>�*W���QB��NM���V����/g����χ�l�n�gA�-��v��~!�L�?O9b"� 
���n�p�JB~��E	���{屩� �(�$J�.�#�������&Q��e�,�U�-Zg�V�S*���n8������{��13��F~��6f�(�S�#n)�åSf"5�ʜ��1����c�X^�"�{A�"ɓ�;�=gc����8������q���'���O�H�*���݉ʜ����0�4�ӎ�=�s\�;9ŗ�;����K��;�5���Kq�E��m.�p(^'���	�U8Xu����?'���Ջ�BB�m���J�N�t�C�����v�I;w�#��{��xǏ�2�C"��$I�֍5!:U���n���JL�.?I�F����;x�Z���z���!6�ڧ��� �osZ��%��јz�?Da6�$̍����&���7o�rRwF�hI���+_��6{����d&nx��پ$)e�K@�TcR=F�_�ȟcX��j�S����NN)��.�B����h�N{�	 Ȃ�����FD�p�c��yO]~R_n67�=A�i\�g��F.�;�[Յ-i����Wn�ؚ��t;���݈s��=ِ����i��I�Ǳ�Zn��/��p��;"�(#Tfˢ�e�-���a�� �����{�o	\a�4�?p��k���-�zaѯ��y�̞�L'�m�(
w��q)l��o6D+0�	m�sS�}.Q32.�s�<�oyY����2r�H<]`I���ǾY5i��j:�j4B"��F�݀:��F�li��,x��=�Y�}U�%q`�u�j&�.�07�hpR���%���	�(���e���ݏ��[�z՝I�&�P�L��z���P'�CeVPDr��"l�}~��QS0�kR�wC���|f?tƏ�<����*��N�Yē�g)���o���y2}r��XiǾ����bm�n�.��!h@�g�v���u�
��>��o�^��ۯ�s�������73��Z�T/��)򐘴�I\���Q���;�m���]���.DJIS���0	:N�^)a������,p��Hh�"�v�c-�%L�CӚ�����OxK-l�0�J�~^��Ym��x�U]A�fr5H�OZ��0�݉�	2Y�m��4���pD1H��rU8��|��^ò�H'V{!:��ܺ�Q"±K���`��n�%TE8`�T�@������)�ƕ����E���s6|Unk3dǧpSG�0j�w��]����)�/�[�y1�����6yE�R�Qk�.�2fM���;��-K��iWq
<�Hl"M��iߤto��"�i�:ؽс�����[�m)��鶶�����������$Һ�xZ��Z�ʠ��D���Aϗ��;�p<�<���t���n�ك�x4 i�D�-��Σ�]�έO)yd��m��9Bcc�q��JD�eɛ��$�k���6�H��0O���o��[]��������z�B�6S��t]��a�����Td�G�/�7��˽��n��ˮܮ�ëoG�{i�����8	���J�Q���b���R��!���r�]Opͩi�fv�-x����8(,��E%ͤ�h�\"��>�t�����.��}���#Zk:���E'm�,jqu>�S\�c�&�v��k��k��/�w����%*�_3]�4��(���%�k�5��/8�<�(������RY~5�E}�C/_
r8��.�����j��#l��Iǹ�$1���83��h&
B������eLd*fj,;�����n��5�wp9H������&�7�R1�����B��8Tsg�m�q��"n�m�b���'��f�M���Q��k�B�/�/��^=X��B��ni��u ���wuR_���MA�{0M��_�����*:�~�$��8�&���������#�ȶ1��/9�`�Tw��T�+2�Г�=�ښ;c�8',�H"�.��ꆸ<���Jg>�֖��nR�[�GP�m(Q�d���Sri{�b"_Z�uN�pO�a��X��BC{���6o���Mh}`p9![_qM����f�1�_r�����e�u���?E	���h���L�c�Ds�(p|Y��t�hd�Fj&�{8��!!���2y.��>�g���G�4O-Ԧ��ɶ:�F!�^���Ԥ�q����1�9I��U5����P�j}i�+��kS�q
Z��e��MÁ�����;�|�0�R��kŘ�1��{$�N�Iz�ǋ�g���|���������@0U�W������@H��뮣7���/\��Ǧ��W�R��ɭ�<)A��'�<� ���"C�T�*�X0�s�:iq�UP��s�;LY�(��� x0�A��Y�.�c�
�y�(�0x���ر�%�?��9�UV���>�>1Z0������d%a␕yR&�Tp7"�����˄C.�@��ƒ�>��iE��$e	�hfϚE�\}5��^������f�d�ϟ��_��3��;������\v2N��g�ե�^0K	l7K��p��
\���s(v�-��\�v�4�VrEۼ�c}��Aus|���HX�f<N�N��}v%�`B�	�턶;�<|��ߤ���bɕ&�5#��9�`�"龾>�6�3���������7�G��!'t���Z�y��t&��|�I'}�����<�H.�4fEX<s�s'�b�'U�>�',T)-��O4���]�Y|}S��b��ƣAu1K�s/����pA�"�J�*t��T�fM �>�@km��Y\|���Ɉu2:�n����u<���Of-�`�B���^Gk����]��?e�=���S�E�y*Pj.,�{�ڔ]�`�I�LN����_I�C�)$f�L��5�/M9�F��y����Qz�x�"�}���]5���k]�A���v��h�1����q������As}p�tj��^xa]��wt�{z�B�ޱ�wܽ�~��tMr�, ��f��s��:MJG��c��PEH2o�%iA��� �
6�_$�5 �m��`��%�s� (�����K�eY��m��L	�ʹT�[J�f ~�����QA ���=�LV��0;M���͹$?6��.ϲGK�˥I[˾D��2� ,Ϥ �mԹ��Q��3gҊ���_N�?i~z��ܷ߾��!k:kR���2}g�q�*���}뭷v &�F̺d��2ӋID)�}_�]9�oY'aP�>0]%��6R>{�MF=����0�M����*'S�x����d��Bf^ˣa�!i�Xʥ}��z�<�v@�,��1�MU:%����n���4AN �t�uN�6����SOәg�I��Ƃ���o?�"f��d�?��U`�!����mY!<���,�,��p�S�2�l�����t�C�ԙ0==ݜ��2 i�l�+b���BEl��Ծ(k�e�f
0e�pe�U�����!a�����)ͺ٪<Mڝptd�* P�j�[߂���Ҭ�� M���R�X��N��9�����P���$���?��	2�/��S�}ꞯ/�z���ĬY��$A`=[��>� �`��fp����|��6BN�HP��KH��s����m��A<7Q=%�2�or�W4KҞ/"n�\&l�ls'�7���Q���6N����h�5�9ڴ6��m��smD�'t�D����U�h�HD2�yOO/Ӓq/b�	M4mɁ4�q����9�S�f(��Y�
E�?˯�H�-��#t�9�Е�.J�2�g�dj�����v[��w�����4��d[�1�&׹�j�}a<���p�Kh�� `��Ǌ[z,�/�4��#�ҵ/*�y������D���*���ZgkΘ�f � mY������#�iI�A�(kj���
���JF��=��퓗Ӝ�z{i���t���t��N�%O,=n��}�;���h�y4�l��L��oL������z�)�c�=�_L�;�.YL�wL�&��#\p���������sQ2�h��	���}�}��)��V� ���y����F���[8F%�}�7��������X:�pyB�4o�ۿt?�D�\W� ���(͈h�����V�Ux=l�VX��/��p<y/Mb��o2���s6���7�L_�җΠw|���Z8�NOi�$��2��{�7���?Nw�q��>�� ��-���M �'��fX��@=fE�@<�P�-�Ԭ�2 ^M���R�}�I<�`dfgv�c�I~���qcY�&w�M��.��彠D�?�j��N��!w�M�7�������f����*��ؾm��:mz<Va��e�]衇���G4�O�����'.XY��D�MQq��Sˉ 2m��"�d���g5��^`��d�M�q�$M�g8ِ�N]�Kp� L=dI�F�T�O���/F��k�j�Rb.�aH��׸�PX��*�9Zh��Qr0�:3//��x6m�TF8n�xl�~8�Z鲁[͎�l/;>֣i�\6y�k�~D�-���|���r��`�0$�O���:��,!F��rvoqh\���k��T=nG�r	����TX�x3�>z�@?���Ē����~�����Gn^��G����]ʛ�MX� S2���o���vӔ��GK�Zb�(��ɉ��vֳ��,�N"�a�3��+�_��%bl50�k`�$���j��ŀ..-�L�ڗ�*7��M��e�<R7w��0b�������C��N�gY�aH�H�5��E�D8��04UM��`�6�`49\��t�Ygӵ�]�����
ޫn�f�&�dv�Wp��9$��E\�s�Zp�Xח�N�L1��������
#�c��6�3/�	W0S= L4y~i���9��2UNf�����T6��7�'������%�ş��x  C`e��o�<m!ʅ0��tQ��G�j���0s�q?��z��"&� `�- d��=���t�׿N���t�]w�husR�T'
���7>��Oъ+D�Ҝ��*�!K�=`y�V��Ub�; ܒ�V/t�T�K<b��H��EC`�l{�P�c�f��x��Ǹ7oB�f��	�� �QE�䱞�
�R���|�0�(�h�k$��&�a��c�I� o���@�6��]��_��sfˊ^���.;�&��G��S���e˖������e�ӟXU  �iem��I�I[le]���<`e���4PaK�J�"�w�J��l2�JҌM�t�l7���8�c��:�K������=��L��z,��x���捔sY�u����q�l��U�KSy�,��(IQ%���}��ySr ��� 򳁨�ܸP� �l��>"��M+ae��K�����a, 480����E��g?�)}�+������M���x2�����W��n����sO.�W�p��.M�Ò�&��S�5��\z�����m�d�h��y�rν ���~�E��VX5��`*[[K'Wj���#�k�<�!e�in�,���s�Z�M͢l����� �$���)��p�=�A����н��e���o�~z���C��	?��G���47\D���]_�pa�<�b�,�Βڤ�Պ������	}��=�ŕ�FW�g��9v.��D`���(�Df��)���*��� ��ϼR֝8����dh���Y]]ۦû�m���43��W��D��ΖY��<&=�ē��������Kҝ��aB͸08�]�?������~��BЊ�y�^B�����^'�Ⱥ�D��֘���" Ȉ��m�XC��rq��&2���U���cp������eۭ<��*�X��p!!��B���� .�a�`��"!3L|QЙ��
3U鑀���IcT�l3�E<-�Y�ı���n�d���9��#��믧��ڋ���?��9���_�M�㜚�A�n��4���?{3]��^!� �Dҟ�;�X~��������5��֯�&\k�[��Ox�U�!l�rN!%&?�s6Z�?���o.f���)����:��`럗}G���6�k�oF�6�w��ų�	��������4{�J�HYAz*��:e{29e)MoP�߲�$��֤�����7�Mw�^�/q}��sӏy$>־Ymy��l�d����U�yUr���%<��Ϥc]�lF�e�)'�`�m��L2sq����0�O�a|[��VP	 i0�z�Jҋ���e;k�r�eB���&���AzK��� Q�H�l�B�ň���iz�5Ƨ�:��γ�P�+�l����qJ4���U]lz�'}�n�������;,�c�4�l\���8� ̑�Q�a�02.����"D��If��d��h� ����ki�5f�(�(K�dȿ��Z��Z0M[�?Ze�U61��� �f��͌�L�L��}�/ � �̢kn'���L�8��s���C�$�#l�m�̈́x��i���K�y��{�I��{o(��i4�8��2�������t��L ���$V�N�s#��}���\���rhʵ�z2����0j59Ӳ�Ƚ(� ���TV�d6��|��`������*L�8��*�����n���C~g�������:�,�e�r&������O=�ԡ/}�K4}�tx�F�*�P���28Ч�^o��US���n\ڞ��{A�<@E4J3N�=� ����4��1�` pi����X���U�m��������z��6�A*�:X�\k�x5<`��a2e-�eB��Y��YI6~�0�*%X'7?��c��cƮ����Z��:�(�w �h�i��x���.��G?� �8Bd�|̭�G���D���<L��zM�r�P�/������7�d�� 8�" ��+�f���xl�7�\L���ʶ�8�ybԿH�?�<�瀌|&�"=�����M�U�܌e�!����V��i�k��g�ؚfΜ���s=��C�m�f�4l��L�#�<2�0��O?M{�7��p�r�0ڥ6m�,��T5�# @7;n6�I��m5Ÿ�}�v���%f -��Ń�CC�hf���b�g�|G�lCCe]�,�"��ؚ��Wy�b[H�����G*Y�N��hPSâ�6/*�uj�#)��P��X�N�i�Z4TE��� �c�/�c>�	�#�3��qn�d����oҵ�^K;�3���\�'É�$f{���<K]F���  ���R6�B�ێ����=�֫�v��Zd�!�HT9��*�b-v*6��af�ٕQ�k�YOˠ=@w���w��� :�M*�L�K'�L�^�y���g���(�g���Z:닧4����qMG�� ���/?�5o�<~�A]ec`�(��Hb{¤���qe�9�A�u�Ȅ��dV&�V�2'�f"۝$�lԻ4�#��\�q��4je�C��0m�P�?�r�ų�|�\ƻ��=^�뒽.� ��7�񜌝-ǣe9���l���M�c��*��Ui�؝y*܆�B�2��Ny�gBi�Ga&έ��`��l��A:�S��{�4�Ͽ�Gwݕ�q�e��ǝm��=�\=��0�RL��ً�f@�'�*,����g�o8�ȳ�����e���ʩF������p2	}��.x` QYe�U�{�LR�����>Ƣ2����WZ8�b7>�Z?3�M�4ϴ�
$%`�o	�����/4�$31���A$��8J��6�`��˝{��z*]��s�='�*�(2�����؞��0M��a0�,d�L�[*��+.cY� ���I�8��ņ��N�KcKKFy=�#���s)-?��g����9������d\�( �(�kY7\�KL�6m�g5���	.J#(�8d����f̒%����x|_��E�VSh�vs�ʫ������������<h6�ӑG�-W���e|f�|��o~�YM�@W��~���#�%�q�/�1��H�K8���{hX1L<���$Dֲ�KW6@Ӵ�}-����"��1#�W��mUXkb�
�.Cթ�w�f=1c�6C�8�鑦ef�A(?V��4��Mq��]}S�\4�:�}�V��ξf��>]q��y=�a���@o�@��Vi޼y�._��fϞ-ŏVb,2�vI59FVOa2h�q�m�+cQ�R}�\�{�ѝ��tpڴ%�e�PR�9l�M�v����6t6m���o����$�� z]s0�}^���3߆�`�6��Ј���^3�7�ߺW�J���P�"��%Zw�%<ư /�d��˔�c���P�dfm�-�����f<�fK�_}���{��hڴi��9TFiV��3���dP`�J} �pG* �P���6wل����A688D�W���%�L�{3;D$��`��re�UV6LZݖ�Yc4��x~&=��g�=@�<������`��\=F�m��؋x<�n��QzbM��������~v����Q��K&o�y�Gފ��Ƕ�j���S+����( �����g5(}\e	�L���m��+]0j٪}�����I�%Ŗ����'�ԏ���*��lZh	�q� ������N�AFj�.���QW�Ug�V�@v��xg�
��0>�3�=g6=��#tƙߠ%˖�;|�;5��ղy���o�ۋ.���c�=���j�Lr1�UR�Cp�۠��~�"� OFCdA���C��pP���"h5����[�j���*�lm��� +.�'c�gB��t� 7M�sĦa��(���c&��:ެC;�CB�hΩH]���M(��w��4�<�s�'b��쓂&��M	2�(]��C��s'�����(���7AG�	��F@ �V�4e���YX�>1�.iJFփ��@���L�a���{�۞9���.�x�#��*��SR:o���$�e���x�����2����lXm[2J���:X����X���6R�Dy2X����Yy���=��z�u�B�\7�5P����@�M��f�\���Jg�-���
�	16�&4d&ɐܜ5k�ѐ.��%t�]�����z��	]�P����f�M	2��cʙg�IW\q����W��X�8������"�M��BD0���o�Q!�ϞK=��ܿH�X�H�b�XH�"N�yT�UVYe���	V&��h [�9�[�%��1N5��Җ<��&�#[��g�0�m��I��"�z�X��1P�qp��eܲ��;�E��qG�ܫ�l��@�UC��߮<���We`���ԯp��g�8aU٤��t2�Ӯ�n+��DZ*ES��o
UY�.�(�dP*�W%���ge�U6�M�Ƌ��s2�� ldD�
��K)ƺ����e�������-���f��v�iS�w7�@���;�ϯ��''�``�
d�K���В%Kh�=���-_����@�L����H��H>A5�̊�^�9��Ȃ̃����e�����LS�w�4A��Ye�UVن�v�l��̓��z3�<��%�0L�h�t�����O��$�;n���.�{�zi��f��;�����^��2��mS�Lr��������;��O&��S�9��d�#�K˚04z�E����Z3@������oZO����,�T e���_��F���cu|Ƿ�)�خ�� {]n��3�%�q��r�L�3��v,�kƲ/�T����*`�v�9s&�v�m�p�Bb:��vo�eo֖ �
d�o|����Ӝ9s2�K��9P�่X����[.� ���^�=L}�����$}*냂2TOً���o�qS����n�{�d���*���u��!�2OFZL��~6!���0(Ό�8�(Ma}M)�Huj00<Du[/�����sɥ���9�U��M�.ۼ��M2U��?��`�x�E����d�y�0Pxd�9�bNr0hB7�V�T��16i�<�Q��l`;�Hs�	/'�L�~5�ݶ�~:�}��g����'�N��#���^�ά�0�� _`o����~��Fa$���R��i[ h���}����~:�߼X�l�M2�M��	����˴�$��H�%���{/V&�օk���\��c�0kB1K�I�T��N��C=��t�����*[_5wir���0/��t�Is��55���qp�?_Q_��~�!�#e	h�w�m��2x���麣�n��S6�`�@&�d���?L�=�Xۑ2����	��S�႞��r�n�nf���F�j�u��*i����0�ZI��b`��Hc&Y99��%�>.�AA[��5��7O`]g^�_�x�-���d������a��*?�	,�b^��H��sȵ�0fb\L��f��8��*%f`��o�(��Y&.���BM��Q��n�9t�7ҙf����3�
dT6H�y��u��\��c�R��h�2�
ʡ���&d���Y�O�K�L�'�Cc�DTMUL�O-e9��*����m*�4��(���iZG���|A^2c�ʜe�0��B�Ye�m�Z<�*ϵ��t�M�ȣ�w;x�-��V�&����~��_�5�\�*�
�*�+0�MȠ���笨�_֤�%5� �&BeT�rC!x1M�������0e�I'�.r�F�Ή�w��F�3�=�ɾ��y6�Xe_��Zh�qAF�'�H�wwQ��!
�x��.L�<��o&�f�[c@�(Ό�3Xm����6:e�6����,Y���#�k����.y��К��?��ho�/Z���"��xd�#�DuO9�ƹq�����6�y[���������h"��`ø(��ӕ7e��G"gn��|4&�Q�ɑ���0�$)�����Σ�x���f�͌���r��Ŵ�6�d�`�D�±{1��pe?��:ӑà��d���f]*d��A.%�z�D�+��E���r�VK�[Qf��>�9���f_��T�ֶ�~:���Dg��t>�J@�M�j�J��IDo�	�e⚺�x5H�5j���0�8lQd�K��gT���!�0u�TZ�|9��W�*2��5�k62m��e�q��d��+'�D/LZG�H�Chҷ5.��J��Ɩ��ʴ�%���DCmQV6Yd���S�gTսTVYe��ܰ��" �l��"���Dt0�F 8u`�D���]4�ҨA���f��3�����{}��f�d,X�~�_�Y�fQ/�����u&�R��Hb+���W�ދ�aB2q��,����p�J��dL%�Ie����
h*���7�$c���J{�@���0n�������#5�r�*/7e��bN�� 3��ڨ̉m����ͬ�_M�<�0�~��D�U���6i�F��47\D���������K�=���N�V^H���p�.��]�ȂS��d��d �����4+��P��f˞�Ȣ{���
`*����jy�^�N��j��
��%�\�рDT�r�f���9�$��� ��>�	��� ��������û-���X�iNd� ��b�.j���X �YKV�a*	O㖈�&iL�Yf_2>��@
1ؠ�L��=)HAH⚬`U���Sc��0�,+]����&g���=�=Y�4c�˫���(9�-,���l}s1��x���O��]���_��R�r�o�w&��~6� ����[ZC��S���IZ��8ɺf��3�AhJ�Ĝ���c��&6��Q6ޥ��`2n�F����3��~O��ͥ��$��=t�c�:�X�L����Og�@h2K�$��%��W�|�y����8�������37ZQV��3��*����6�[)K	���Q�g<�NC'=�I ��P���Y�̾��Y�9�5��ј�!��n��X�;�E��&� y��Xz55's�-�4��ַ�����#coÂ� �_03�I��.�H��������d�Qf�'� ��*\����*�h�.��Gj'��I|�����<sWM��f�c��zʟ5A����n(�0 ��m	Bm=�=<�^�����V�{޽�G��]�zt�؎�d�>�(�w��#��)�x2�z�Z>��5J�K<ܜL &N�FU�5�/���j׸�t�8[F��	�K�^�W@c��'�Y��s}�p��D
�Ǉ���_����ZJ�<w�O���[`�X�Lۏg���4ʢ׾�N��oכ�n��1C4Gyl���4�l�Z��K6��k�uM��5=��3�_�?�#n���/���o��w�%�l,��-Z4��������=��w�$��՜�U��D�, ���u�8É��s1Ъ�q[�Vk�;]F�*��('��T<�y�_��O]şqhm����hbՅ���?X��V�<�c �D���ڷ]���߰(��1S�*��t%���S�b s�˶���!@�H�ܽ��<0u���@�]eͽƽ������k�b�?��hy��:��4��n���6��D"i6h�Mn:��'��Ƴ�v�F�D8!xY0�رRm��s'2>r���Р�?BQ:ա��k�q26��2d�P/�\��fȶN��V�?�� �ēu^�Wѝw�MK.��?v :{��o��ݻ�͔CgX7��@&���iժU��ڱ����܂ċ]8KքA��1��z1"믃�c )��㬪?�u�d��%��ͅ5e�)L�X��2�C�dߵ�p��^�����߇k�k�7.'V�Y�k���k��xX߳�>k 6Z�>��5�	 _�A�{q�Jk�󓖭������G���U��̍&_�tS|�[_�5��d��5��ʕ+ĦN���_���xT���?�
�IR�do�EO��j�L?׮���W#8x�|��,�z�N��R�+���6�E��Q�e�G{�~�ӟ�A���@�:bs��Gced��������h��nn�^b�4%�4ϗ��u���r`q8�:��<��i�\L+je��r��\��YҘ�kq'i)���
"���܊�h���C:����)����$˕�H9A\�իi~��~09���ږkL�3� ����5 f������h���ܽ4l@�����m�め��_�x3��B~�X&yO������< ]j���X��ٳh��݇fϚM/zы仾WX�g]$ 
&	���1��_��1�3i��z~?��6!�|6���ؓ�M"���v�{����L ���٣�Bh[�׸�&&�ͦy�؊1	��s4i\�q45C�<P��������]t��c�g�> �9�|7�p������\$ TNl�&���Pty��ϙ֙���bq�#.���ƖS'���Ѥ�^���y����b��v�y'���������5W/b�#x�����Y�0���u�m�]i��v�_0 ��@����[i��H��(جɰ����N;�>{���:X�\�Ȁ2ER�:n�\�=� �w�}|<f̜I�ke-1���痯���nK/������m�e��ܓ^��WӞ/~1m;s�|W�a��ϮZI����<B��?_?X�_�=��)�LkA��SP��R3�xl�*nu�����qOs3��M����"u�f�Ci�ȑ�-D-:*LN���f�4h&	�=�-�o���ҴFG.�}^/Of.�ѢգKϹf��?~�63��ló��֮���]>����*�� �p�4�_�6 ct	L��ny᷋	_��o�Y�H�4F�ُ�٬��H�0�8!f* �|ˁt��'���3��?t�a�~a<Js�6��w�5,���[�����M�y����׿�0_l��V�:.��2��O,y����������M������su7$4�.�Zg��=�Fx=����p���+��#����|^Gr:��>8䒒T�����s���2m�4����7��-�w���N;��E7��-��s=��9e+���㶳���{��a�q.��]|��t������1�98D��0mk@�����3������HY�K����W˼����%�B�����G6��ά�h��h-Do��ē|^a�a���!���I$�~t�D_�jD�ӐҘ���dR0���	.y�%��Ŵ��5����R�{�䟇�=h�z	�g~x9�<I��&���ҴsC��D��zںodH�̧?�3҇~��o?�x�[�l���2��
��ijy��6�����htk�e����7� �9L8 ��k�8������u �Q��f�ܚ���Bj �:" ""(��H��� AQ���NPTP�j ����!	!�BInHrSn�6����sf���ۓ����;;;�������'<�ЛI,>P�q��9��T���	�X�@[�׾��P`���w蚫��;３��XL� nBX����^��:��TsE1?�4�b͋(Ec)ff��L+��X	�	�:g `�g\Ig��67��0�_o��Z֬Y�|5mџ��Ӝ���qFt��h�ʕ4b�H��|@�JQ"��PCM�� xʐl���~�eL?c�T��rIg�~&�r1���R*v�WR�C`�!���V�R�o̘�}��s�7W���ϟO���T����(�V]�dP�,�E.(�=1��R��\?2�~����w������V��}���ӱ�����rꩧ��=�jkkH�3���"�O�gd�/"6suxb_i��Pc$Nu��t�E��ҡt�-��?��j]���F���#F02ms�|xx���I��q&�L������ŢA�GJ<�QV��}��dę��%b<i���XO�V�K@��UB�<�ؿ������Ы���g��<��3Y�w[*�4�L��24Y=U�-6���.�򢻾�*�;]�6i?�c&��yN�)�F���#Y���e��/�t���WO�W_z���S\���$���$R)�V�*��_S�=xx:�iS 7��]�o�W��`|�V/�y$��ޡ1���7 ��v�z�t�P0�|��s4���%;�3\jI�λ�g��$QK�M�[
w���<�=�?���t��3iɲx.	��\:�72��FLEc)�X&#[�@�D����J1X���M3��Ъ��_K���@,��7���3���JFb��~����P�	,Ϯd'C�)�r��̨���9�d�LU�#�4/N��q���NHj���dTR��ղ5䔋zw�gK7<�������S�����t�����T�yO��1.�k����l��4�ι �#iMGTb3��������WE�l�+�(4,Q��y�9^B��kC�U��~W���Ǌ�CLL�n��,��K*-��t"d�qW��;�|9S)!����Ju�j�2��9�[t�i���)����؞�5E0�,0�:�+rd�]4����d�YK��=ƌb��H���Eo�搣%<aV�@�}6G8�)wtw��s� ;;;d_�MH�F����dt����ʌ�%�eV�. �|���á3.Jsˑ��:���@/A�.��w�MO�:!u��i�[��z�d��hã�>�	�q'��XJ*�� �'���֩�h�L�٘#�����2Y���5k	[Z��m��T�]R�k�� 2�Ѱx-}���i��WhŊ�4~�i]��k[*�R٢ {[p�LƏ��ۓ��/Ǔ�d֢�+�y\3�V*9ã��Q��D*A5�x�\�.J2-v���X������a�F�V�Z͈K,.���qZ�]��1���f�����C?CѠeC���.�ݮ���]��{|-Q����U ��� ��wމRu�T���`�+�E��pչ�30�t��h��t���G��ռ�z�T���@��옩
c3@�I*-G�[Yhy����Ķ����}X��ce�R����;�C�������qN�G��:�[4b�(�.cp3������l_�rQ��b��O�)���0�)\�x�Ҫ��[���*Y�V�J��	E%��W�]��'�es�G��s��C���i℉�_����� '��s�~/[��p])��zF���7��*H�����kx�b�B��_�HS��W�����{�~�qz��ghXcS���|�ƕ|������9>�䓜��rҖ�o]�*��]]���{�e�\J�~�	g�DY0����\#鵅�w�~��`�Rjo�0ژg��e�E����;��8�H�n��(nE�ʬ��@�5�<��J���V�ۧ=��?�|��_������ι�"E���ĸ-rv�������F1jW��@5���j(�s��^��P_�J&�.qeC3����>�m�F�Y��R%���Y�����F���b8X'Т��(A��ȓP��B�8����0����y-�y��S�\1=�R� TPC��SA�(����6w6}�_�b�f���~���He�,�Û��:�U#�,-<��q��V�,�]wٕ�>�h���,�q����+h�G�F��Q ���sw�3��e+��CRZ�5�K@~�b���@ds>���8��j
]���H�`څAV#��@]��h���{�����F}��G�Zx.�Dվ�d+ќ��@�̀�	�G�ʕ��PƏ=�8m��t�����e� ��L���bG���x��:�4z��E�Y�a=/������/�F��K�9S�g��m�%�/�Pm�7�V���7#�>�ўy�Hz��閟�|��7�WG��_��2*U2<m,X��m�6^C.���d`Q2��+#ٶN�ڤBd2L�Ā׶dU�%]}<���
/�NQ����x����1j��p��v�*�z�P�Lo���2-ٜ��k./
��q�
��ʦ�CuDz
�Q+��w�=O���ъ�)��^�^��Fo*z\�x3�Ĭ,M�eKO�a<R6Wࣜ<Ϸ��Q ����zr�!n�U��������G~ѯ4�d���«���k��~����}통~���:�,�[��A[WS���z|��L[*)�k#���Z��ۜ���������5
�OF��Y�{�m�滋i�̛XA,|�e���i��1�[�󍺸?H]x���P�m����s���<����"��i��i����&�%������.�%�5r�V�]A�a
�S��!ڗ��D��\���mx���#�
�w$%)�\F�e�[�팣�@�gG+�'M�66sT� ѫZZ��7�.�"� ��ZRɨ$?�ワ�[o�Ŗ�#TKJfc"��^;L�i�����g��j�8��R���z1�%��*�9Ʀ��o_:��S誫G��ײ%U��@�G��¯��J��9�����:���]��c�3�fH�m����%���W�C����*��eQb�]<$�����H������Wαឺ�O�O{��p��駟�^Fc���F��kx/0}C�����24�����?��{꟏���+i]�Z.*����d���[xj�����5r��Wћ���3`O��	�s����m��H���[���L��a3b�5��~vv�o�I���6����
&0��kiiy�.���@1�|�'�y�t,�d��=c4���N*�8*��LUɔm�����wvtS]}�{����hֽ�0m�+��N��G����Bs���6B_�ET.nCV�����EZ*���)�4�1��e@�m�z�]�b�n����:KZ�y�S���> �O�z��Wy.�bӨ\��k��l����q�sQ���x���k�i�P���-��
�9�O8�w	X�y����N�g_x�n��:��hn�J&Le՗g��r-鴏4c�Ɩe	�
�i/��،#C��.�8k*��S��:(����K�P3Pn��M=�~�ᇻ ^�"��2J�\��ŬZe�����0'U�Y��'�{�x�5Z��,�ʓS�3�Dʃ~�
k��Ϧߦ�B٬Sd��H�bO7��k3��6�e��{�<���P��S2�xR����B�*�<�=x�_���ӧ���O�6����
f�[�8<��um���3
/`P�HAX���	U:��e�����_��t��ɓ_B�`�=f�m�X�J`++�jDJ�sa�dk�zQH3�����l�"�rp�4��9��,�5Ǿ}�����~\���9�2�c	�4'�����-ZD��Ͳ ��Ln�0�Y��6M�e�eX|�GI?l�Iܓ�Z`��ȸy7��k`w�ᚡ���p]Qn�ɼFi�_�����w���`�X���X�=wߕ����rZ��B]�⬯�����ù��u)8r,���??�¢'/P�$���.��b��r�'ƭn�_OY���U�x��NeϠ�^\Us䩿m;���=��aM�d�^h��ko����p��݌�ݡz���쪫��7�|���z�ytuw���E��'�P��#x���Ψ1c�W^�뮻�>)�L]̡��3��EL"�:�	׋kt�q��Z2��L[������t��V��u t���hM�C��n���aR�e��"�)C�&���m#gy8"���R}2+W��D%�МZ0.�҅A�6,�`d9��m���˸/�G�Y����b_�(dDB@m.�Z9��M������|�9�~6Ҵ�;�EK69�!hl����@Ͻ���׿�0#��=5h� (=e���2E��ϓrdŊ��P��/}���U���T �P<�����̳�����d���_����x�:bG�7��t2R��ܗ��Ҍ3h���� W@��Ⴠ\���z��4����H�>,���L&�Z#�MY���Uh�T>9�(��?4c�J�'�!���Y'���5����x���6��d:���|��`�N^����1V>��-kdC)�U����daĠ��];�"�|�^���(�RF�7�t��Ri�����\z�W��w�!3$@.婫�ηϡ>z���uu�3;r�ϣos2��</x>CBh;��2�1��$�8fJ��-:Ղd���V6�>��O��R�v�ܿ��r�5�n���S-�AS�s�C��#�5�aN,'�s�﮹�����v��-K},B]b>/_����_X�[2�EX�R�̈b^6���+�H�a�Y� H�G���y�c���?��������}�є�dx��$�����0���W��|\vn�ي���DU32�� ��d�����}�S*�U�bz.ᔶ\=j4���`�P4��~����>|V<��~L�f[��Eߣo�yS�5u}���7�hm���)��n�Ȃs�A�6S&<���cBZ<?��C�ҲBv�D� ��J�ýg6*���y�'[x�
tX���SOҼE�i�����~3���Ř]�!�n�/T%+���o�s�F�*��r��p�JF<Ri�I�4j�̬���~�#!"���Q�xL!t����Gp�E?�Q�.��W�L�*_`[u��<��2�'퉰�%A���t�Umr0v��=���\��= ̂l�f����sXٗ8ΰq�K� � �-S]�N�z��q�Զa�p�u�Ͼ{����&��vA��=����8����o�ʮn��W/�T,���V�h/�)#q>R��R��"��M(���F�I'���u]��M����Ѻ�.���[�S]F�]�b
�������	0b��^x��\z�e4}�tf�~I3hj���.V�DdKa4��H@�bۘ$|�zj���萙���MU�i��AY໎�w������j��wt�M����E����+��wev��s�e�Wm�����U2��{�-��Hfd��*T&k%Q`g+�^��
,p?!��}h�B'��m������FRY S���s�*����/�8?�'���wd	�1_�"�y�]�	JnvGW�dmG!1�p���J)Ag��۞�Lي:�"��3�^(�c06<��c<���O�����J�,�N��ѣGI��D���oz��� � �"b1C���a]s��69��@�6�]��y#�
P���	�Z�@��vZ��.�w���,�'�92���w�D��иq��I�����nT�J&��XX�
Cp��YӲ�	c;")b,����Ν�nX+N��[+��э�܌�>��=w#S2��p��GbN_(Y���({57ΜI�Ǎ�SN=��v����8A�(��4M?�n��:���h���e���Rn��f0�1�;��,]�A!a�[45��Owu�"=e�d�J&��K��T��E��eE7(�}�Q���b��.1�wH'<n��Jr�M��4r�>��=P;H�[��p�TK��L�����AU�����ba�r��tѢ`�0,�ft0�����g�3�>K/�������޷��=�r�L�7��p�;�@]l��|���y���E��w���TG��Xf;Q"�ԒZ�

F_�[������2�Ë�ࢻ�����B�&Of% n�D���QƄ�9m�4����_��K�Ҥ������RE���"\�͈"�R�$Ղ=C��L�
�Khȋ����f�\+�7�I�����!�-`���բ�q���5�TU�/�7�Vd�i�ʬEW�k��=�k�2ƾ�}�@M��������������#'C���:���LKKK��#�䁡9� Q#	E�o���h�eY�����W�� �!��~���֘��J����4s��=���,��J
/���7ޤ��gt�n񿟎�$r)"��v�����Bl���u�xaq�����*w�қ���39f�����Qyw�R�H��ët�]���54^(����W�;V��ّ�p�S���Qf�I�J%�u��جy�!���7e��i��^�Nn0��ؓ�=?̥Qf�����T��!�I_�k7Io���R)^�����d]vY�P6�a����R2�
�	��~fK��@@;�BQ�LR/q�QE�a+d��^z.Ju����#���#�$Q#��g��n�������oJ�e�#-a�H#�މ��|�p�Bz�ɧ��^�ڋѢk1\�cJ!�=�j�D#8amN�<���D#����	���E�x� �S�O���.3]2�Xu��Z��V��}���ϗ.YB/�q��{X�k�K�_������i�ڵl�����	���#��y�=}2����Lw��+��B�Yq��'¨?�rj#@�10�Q܏�x�NY�d)]{��4uڎtо���X`Q{�����ө��J���t�p��R&$5��X�>NM����+���1b$�,S����8��[g��e=���K�G5�3	�I�����29ތ����d2�e"��X�VtR�d�)��'� ]ѫ�x�bJƟ��~@mSuU%�9s�N҃n���y�L:W�T���D<+���3�JN�����ȱ��������v�eg^��`���c�9��~����k�R�P�3@l����Ξ̤I�~�:���+[��Ue�V.$�[�o!	Cv�
{3n�q�l�zD�d��:)G�L����>��s�`��}r���At�3��8����>蠃8L:x4���= \��aY�%�X�"���c�n���(�<If���y���"��\C�["��S'�7�����,��0]Ȫ�	�O��8_6e뭸0��_��.��~w�U~K]���w4g|�����ܓORw���Lݮ�r�n^��ĻV��>ړ�y�[ Y�՜�)�9�8,|7}��/�p�]4\(�� \�}��2�c�6���Y���^��V٣L�L��1����y��fK��7�_3�R�Pθ*���2�S��[3�䃲�s@�!J�4��l� ���!}f�Ԋ�$;�7���ı�bt��R�֢RP��kY�*,��a`�6��uKSF����gL�_^��(� ��W�f�0K����ފ��1.ۃy��quk+�{Ͻ��#>O�=�P�Z���^r饜�Y��29H�hىf��C��A�3�^�����ht]cq7dV�ދ_lI���{�RB"|e���#S�~9��YF���`]�����D󘝨_�W�{�C/��b�9�L��q�d4
�5���醫��V�W/:�S3-�'鹾�Q�e�.�S1Ce��>�Pl�r�*�����>
y �7í�S�v��SO���#LS�M~���U�̄Y&���K�w�4���b����e_�o���X�iP�L+ؾrAԂC�
5�m֏�����qR+�}]}S�<��[���{�~I��	�岹s�2uN�T.|�4�S\<�-@x*�xPq~Y�*&�xB'�������j�F�(5�7�ó���ږ���
q�9ߩ��b��^p͛7��<Sl���_m1QUz @�H1S#��ȅ�X�є�ڜ�c��h�S�=�+�D�g�j	�u7��E��1��h`\�?�>��.�T�c{�(�lɒ%� 5�2$���2FQR��ܶ%_��
v��yx�4����2��x�d�8quv�c��,����y>������\K���4�I�2./�A,VC�P6����4y�m輳��MZ�ʦ,�I\?���bp�}�E6JVx���Q2�����[e�
E�FJ]���
�9�����&�v/�mQπ�$���N$x��?MÆ�V=�;��[��rse��4GQ-��J8'�CQt��f��%@@����,�&R�K��,��^�׮[Ǒ(���{�>���w�y�ϫh�d��QUPeY�������+e�O�o)
&z��`��,;�%��G#F����k����{Lہ�C2�H� =*>�Îtʩ�в���a��jsO�z$u���J	3<�X��4CcCQP��`�I[\�ǎ�Pg��!l�V=Ǎ^4TYV���Z��)���2�N��W%���?#U���hD���a��:�^FI��h��LKKK+15�nX�H�ZF����]���ךy‮j#�T2�2�ʫ/�P��L�$'��\z0⮀�3�<�4]x�w�����������S_>������W3`D3 ?��^AIV0�D�l�S#AE�鈚�}�`0�"�k�p-Ӟ���J:,��8O�<�.|'P�o"��[t�Ǫ�Re�ѡ�k��`��0�u�E؎d�H��E���iFc��?;����\�N$�{7�/��K�zS�L����94�ϔLtÆM�d��l>� ��ʡ�7��f�3���C�d7{1���T�����J��Kl��fFm����F����\���Z:�gаh��'T��l� bL�:����E���ٳi�x�a�1�S�G�A"����o��U���ߺ̧5�k�^x*.����Ph�,���3�^9���:�N�ʗ����ht�.�ή��H�2E������q�=��caV���裏��
o�,����̫d��rA�	tAss��f��K�eo>(XHF�����0�h$P��J-c�W�PZV9���ˑJ-���C߳�����yX&/b`�mT�G>�c�� �L�4ru%�������� �c�]�`���T��o���Z׮��PD���@���v$� �:�Q�s7��"��o��7�ۖ~�ҕC��[?X�"����@^P�����]x(�P�^��㍋˺��SY�$�	�X�w-�5�m:�ﶵu2�TgG;�U�!�2Q�Ǭ���Aߩ���:����ix�)�n��cBZbj�"Cv��n�\����}�:����dқA�0�0L�0�>��}Be�Nʝ�E�H޻	�u�����~E�| ����^�X,"�,sјN*�^�bN����yNY֗ūP�����/�AS=I>��#�������o�2��cx7
�r�PD�<�p��޶��i.���Bu'�I����b�0����!���h}��)�Ou��0��Z�G5n����xѻ�Z��Z�%ga�p�*��lh .�bc���R�R���ݶlf�����ŋy�$�n^��c,d2ė-[`\��R,��L(F؋��d�L���R�d ��g��՜L�K_���h6�{�ؿ��_�K���C�����%�&����cz{�z�g�vF���z5X06M�^M/Ǵn��"�FxA5��+8�o�0�<a�m��9z􀇢�:'W�l|e���K���f�}�}p��۸��,psؔ%P�o�zF9�p���\���qTn4�
��%�Σ�C@	�h�ZZZ�677.Z�`ʫd��醥�G��Ԓ�|�}�8�L��W!#�f����o��y�£���l2�_1��	H;�M7ϼ���n;���O�����MiK&�?�)�r�İ�_h�4t�ev�Y�=��E��4O@��7�����{F��&M��!�U�k8��06��i`	h�:�(�{�N�韠/��������a�X�B�f��^x��L��~�`(��=��;�^H4��s�3S�0�sBo���DK�;�x�&�'����<���{�~pskkk���&e�O�t�4<���.���Q����z	���ţ.�D�U� �E����|m�׶��LS���s
�P%�m��E�ok�l��3g��@�m�/^�����3xą5���;ӗ����'���--�n�z�Ux��3�D��eҖ�V���@���#~r�$�5qjm]K��wp�~y%4�i��'ܟ���?R]C=�k��X�؂��^,~�H��!�Y�����=���M��Z�X55�]wޅ�m�ˮb�(�LSӈ&�g�d�����b���/�Sh�1rZ��FS|���q�k7�����y�Jr��
*���V��������*��M��0�m��
�2�R�mp�x3H6���	�զw�w�_��n��V0	q�#�`VJ�.�9s�����s�z(i�6��J;@��niժ�4�|Z��AÅ1�{�`k�@��_���kl^��q�����!,�;�I�|�c�w�͓F�nb��j��r%�{gw���6;��
 �������q�0���=�Ip`�Ԉ1З��8��	���2P
L�:�s'8��G2ϣ��#̛S���ͪ2��s�K3�Q<���6��c���]�;n�w�y��z�s�9���n��d�����:rŜ|���9��O}�$�1�����Os��/��@ �7�O���[�8q<�r���]��� ��Vww�Ï<L��DV��D{2H�
ǖ�*(�&˜�΁d;m��ںZZ�q;������lأ�@� �x�h�5��u�Lv���Ԗ6S�g
n"�!&��ۣͫ���L ��niqZ�Z�8?sۭ�Ѿ��K3v��O��.�GR&1��{��d���.@�?�.���Z�E�q�0������Y�p�Õ!J<���y���t�P�˖.�[V0��G�ċ=�|�i��u�%��ܶ�f+sk��Y�� ���ާ��z;uvurSD�ۦV�۟��؀7���u�{3]fY�iK�Co�
���ԈGw��Ȟ����g����r��v�O�����z�ba[�d�g�0����!O%J(�4���u3�<I�*�p�u��jlger�Փ~Z�;��ZB#4����}H�����_o�����k�<^�`Xv衴b���QX�PY��e�[N��C�ZLUq>5B���s.��V<q\f�94�̍�\t%DyC���}}�G��~�-XLh��̞�g?����=i���s��q���/ڟ�y�c�9c%7�|�R�LR�utt
���v�c7:���r���gt}#=���t��\u΄��/���[�Z�!����Sj�)u4�N�=0�s�[�KGȖ�C(�������+DgM�h��1�X���z\[>%ԣ�>����s�8��`LzU���{﹧�~�t��vQh�,Ǎ��G>�d�,����1��9�-��n�r;U��5�=��k/t��j�$=��S��_��~z�)
����;%1Wc�=ү��G�;3��7�4�]̊9��)r��b ���y.Ԭa��q����}�>Z���~�	Z��z��D�1�ӓ��G��8�DW���o��vى.��h�)[�ev���g+�|i�<z���}�_�s�a�a��sCf$u�F�q�a�e"p�P���ڭØK�7����Y��-�xW������;g��He�pZ�H�!��������^�� <�v���λ����}�ڋ����g�)�Ż���1cGӦ$�1�e&��ښZ���h뭷��?u �3k�G��V)r��]�N�_��Wt�wΧ��x�ZW��f���Ի
{D&P�m�i�<������!�̬ lL�z��S�=��c����י�ڋgc.�T������P�t*��U��Hbłoe���u�%�� ���_i��x���g	bo8 ��C�.Ј1��SG������א������)�m�����8�>}uc,�����K���Mjn�(�X�6
c��&��a�#�|�b��E�#����i����R��
=�5���Įt�UWѥ����|�IV�T�=z*k�7����|�`��7Π�;���Ɉ��u�Q{�ϼ8�zp��F�
����f<;�.������e:O.�+�,�E�`ʇ'#���7��J��L���A��D.:arhdi��2�oٵ�%崛�!��m��ʎ2��mE�� �Y��]aٸ��Ҙ�sYV������<K�J0ۖ�'�a�U����9OҵW_C?�ɏy��1���iP*�0/�8�h�
,�W��NU� �xY��ph�?C=�߻�#���G�Æ3��o���=�<�wb��LP}M�:�;����?��wލn��&F���?/1sÊ�?`C !����2
�1W��T�!`�n[��(�Ec�lE��v�m7���q�N����|oM̡��z���[4���[Fh"^��<�MT��%d��t�����O�,*c#�f9v(�?Ҵ_��(�u}'��TF���׮]��J����At���20�-k�? �#Ø=_&/P8g�=��E"�7߄��*?���W0�T�ɔ���ZX˖�|���=��;�	_;Am�q-��Ul�������uO�|r��?��>��ϳ+�sl�P0�x�xl����Yg�;G}D{�=1g-[��� ��rld�%�V��q]mm��I[oM���
�=��T�X9����qg������o��9��йmb&���F�z5=I+6f�
� sҒ(Ons�g��{�x��y��_�����:aP�����J���P0x4�^�z�̛������S۲����f���ֈ3�&����_|�=BY��c��v����+��bBշ�ϣ��E;��3cFQc��N�H��A��	f�\��=0�|�s������/�w/����M��"��nq��&i}>#���3ΠSO9�{�Qa̦��x]9�+���%�Ĝ�����9t��G��_�"!����3���c��8��f���o�Uk�PLxZv�Q�w���c*���:�팄.��__[1dr�|��{Y�=,� �K�M̴�+K^�cC�Nh*�{�ٖ�߫�|Vg�i���#��2�F�e��P]W�o��>z�t�A���u�K+���Z9���~�)�R,J��3p�n��Rĥ��l�c���(����"o-%�����-��Z�%K��E^HW\y%�מL�b.+f������ˤ��ţ�@�|�8Z���0g@�ׯ_GBɤ��u�u�c�P[GS�nh�ٝf�X�"�
+ ��-Z�]|�%�ъ���׳q�t3U��O�S��)s��u<P�w8X_�.N��hǬԒ7N���AtP�7��&y�I'��X($eY��)oF�͉#�s3C7��L>��<q����$���\̷_锰X�}C��M_�s[���)KҖ�|aQfč�a�B��f�%�FC׍���I��@Gk�ɧ���o�3�~ʩ>Gx��ʢ��w��q���V�&���ٲK����]@U�t 
��P �������梅��/����9��?*B�+�{�DQ�٠Q�d�!���@h�2���i:e{�R�ˈ��AGW��k������^ҵ�_KK/fz�T9֯�D�>�71�Y:�F�'Q�s��2��R�e"M8ȹ2��҂̀��.�S�o؈�-P:C���
�;�ٹͬ42L�Zf�2����vZ�q@7�E7���AW/��A����'�	��Q|�I�4P4�s����9n��v�sӳ�x��~�*ts,���7M�8�?VJZX��<4��e��F����g���ʏ����&N�Eб(+68B�n�tA'$�P�r�B�` (�@~�w�\C����2���	�qѶ;�٦.:����sIQ�P53�d�*^9���fh���)�S�{�-Z�֧V2P82>�*��	V=C�r��^����':L�j��Z�	O_��d���;hH�� `�W/7o������&.,�7�ϣK.�]{�4vĨ� n�v3N�(�H���&��BVK������So0X��M:�M�ǎ���ޡ���'4o�[t�	_�{�8�|�s�[��e}�d��O���Ĩ@��n�֗��)�(t,U)O�B��=TpW��@���$E�.-X� ����8'"`&[L>1�LV�Oh���P2����1�L��3:S,^R�^KZ!L fB�����/H}��`PXA�u���]w�.;�B�]�=J���s5��@J�R�0*h(9����u c��$o��6W}묳�#���;�@+��XV��@.�~T܆�Ϸ��ֶ�e���GrKv j3��G5��?Q'�-�V���!^� ��v a$�e�d�AY���d\$up0`�ENb�D�J�c}��E�>O�#<��ḵ����Q�Z�Lӳes%5�s�F�B�s0���q�h���}M���&F)u�q%݄j���o��\(��CP�14�2z1����m�ن��ʱ9��±��	��駅�?^%H����*x��~aF@6�ė:�������CA�#
s��a8�Ԥ(՝�����������6u*}�+_aKItJ~-�G]M��R��Ɲl�L]��NaՊ�(&>o��A�?�<=������'���{oV�=���;�*�>�p�/�0<+��-�%mK��&����|�pFHݵR^$.|Y�c�!�t�}h�kx��0(�c����\( ��?�U���-p����x`h��խkب@��#��$�i)jk�k���ʬ{f��ڸ0-Zx����+�6�p���W3�� �|E,�������p�-+��e�Q%"TXD��b�G�"�"0$[�q#�y���q2w����I�&����i�ɓiyKw?ml��tH�3(G���ŋ��os+�z�Z׬�{��
J`���^�2���YU����2m��X�e-5>���i.�i�l�b.�>�¾P�2H=d:::���&�>W�b��^���9��b�\e��l,�_㤪�;�uŢY�n-=<{�X��~����՞,�৫�K��MҋT�X��ǣ=�#F
�%ŴEs�~Z�Xm���w۔�Vr@s+o.���'�A,��]����'/�ɹ q��$֮%�����6�Ae"ↂc��Z�E"��X�w�{�`�BJ������2w��I�}��T2�����G�p6�5J�e�J�-]��\��lqݚ���⻲�oį4���
�I`��J<2V�身�3��8E+�� MJv�3�L��d���t�xϜ\�8���A���x�<Y�D ��S�hGzG�XLt-���T��/��Ō�`Ó�����e؏��ǐYX�` �Ǎ��ԄP뺝a��g��q����V�l|�!����4�i8�W(ҖU�{˖�'���T(�]��׳0���{�}�(����a-��U�?	V�k������j=�(i �H()+��ώ�˗��0�J(���,����F����:�p=�6�s2�{��+�h�r1�U���i���9�ʾo��d�<j"2Ipad�W��K�@u���ډ^H%��x?�=��d+gy�D����ԑ����|�>+Q0��d�x��ޝ�8/ıWPl]�1TB�a4��mc���+��G}��a*7cLD��l[�tT-+.�}M���3sa���!Xt������3�UX���Z��[�cW�!��&a&��=����zF�� �10�?qOb���v���S�a�'}��d����������Z)^�Xt�$�.�e"z^��s!���[)�MU
K��`�����6�t� ���2���M�o�������Yo&/x��}�k���P������I#G�x�&t���^Io�W2��ij3���hik5����4FANT�V�7���|X=T8ds�0�KXr����q�𥏥:.O��!�S�vUyl4����hC!_�L��&��0+��P`�^�ËRDw���-:|%�c��4�< ;`��F7��ń)V�\U���	�-;��F���uMT\J�{�1��<R�L����b^���@�d����TG�������%=0�����^ʠ7�Р��{7�=��'�T�`K��5Z��n�h/�]O-�Jä[Xի:R��Bׯ�	��y$!9܇B� �-�H3A���oE��~�2����5�{2)Bd(����JU�R��T.�(�\�B�X2g�:(aVR����L$�5S�N�����a�[������y�h�����gV�ȥ�
������u���S��q)�r�Ih��ֵ�V���}]-Z��A�uy;�e<� Q����JU�R��#��r�=/�C3E��O��b�u��ՙ�d��%MW�~�C�e]8W�����pv����d���h8v��^w%ŉ�)�ungs1�CW���7�r:���-�B1�JY�+-@��X�7��J��Y��n3E�s!BQ%.h��2n�TY�94'���W��1aDY�9��7CdVu�T�*U�ʐ�<2���e$ƃM栿G:�.�y���!t4U�7sf�n���U�J���e��g��Ȳx��R��m,�
D��/O������m�|����}Z�չ*��B��jN�w�Vs2�����L*�j�P\E���f��?_~�O�j�䁖���7M�"Z��ʦ*P8�*u��N�4�ArG�EL_�^ �&͔=d�y�Z2{��~��_�a�|$�=��7���6�4=�r���h�-*͹��ϗ�ٜ���>��'�3)wܢ 3���*�-���l�P.xp[T��7���v� _+t�~�I�6�i��d�R��TeP�D�iz�0[�O%UF�}�h��Ŷ��e%��d�\��3�R���5ꌙ:q0���y~U��M�D�꠪`�R��T��5{V+n�J�2��4���K��>e�IVY,�P&�X�Ht.�|������{U������JU��dQfd��*�r���]��a�%D'�}�����-�tĎe;e�b��:(�p,~�l�*�f�?�����oF�Y6�?\C�=7� ���yw�u[���V�Z��1z��}�1�R��y�z��R�8����h
ߵ����������[+�7/�D���]��).�#2�}R=��:�f/������_;6��~��,)c��&�?���Mm��,;�\Mӟg ���}ؗу�!ή����U��d�6��JU6wa/E-�~땐1�{YE�.e�߅SgB�c�.��G�o�n�+D�\nZ��Ii�s��Q5�V��I�ugH��`�ٰ�T�.Ӂ�պ\ȉ�����Ƭd�碿l��hr��h�NFa*�B9�j��*CI����Z'S��&f2
�H�KвY<g�6�D�*��Kdq��r�W2�7��� �%�͸dsFb̴��9#�`{ِ��Ҡ%=�lT��c蠜ͅ��ۼ�dKJյT��R�h����%>���+z}�U�?�<����oV4��t�ޛ��S
���2�-+Ó1��S���:�6=q7�����!P"�P��������Rʑ�pY1�z7��FGYn�����*}*�����]�^�^5~'ξ:^5�*W�N���P �����F˼~9��
=�*��+�o�ZOJ�}�/b=N�.�)������z)e�0���2�����sE8VnD\��l�`
uU
RhR��Q%�V5[%н���E7��0�tW�M�R���A���[*�W����M�r�硛}#���V>�m�AY�pK񗱒�������(���z�0{�C.��1 �`�?�kh���B8k�F�ک�2)�+���u�S�r"�`�o����e�y�H��3=�D��ǥ-�<ǉ^��%�I����s�y�%\���~�s1���8E��PRƕ�IbX;�(�-�ub�f!�zrVbU�����GɌNԪ�`��o��:����xJ݁���UX&�XTSS��Fmԉ��[��P�P��[*]���Z���^g�/�<���^0gn��!QP��9����d@'Sr�E�\�V~�e�1��i���ʰ"�y��б�=���/�Ѩѣ(&�;���}ǎP)q��5Ex1]��Ly�2�]{|�f���k����&����vv��9�2�\���DM@,Z���{�Tb�6���xl]���:�(�yn�&{�̅Y�uh��=۞-ԲU<�P}C=����d4��j��$_y��t+/�U��s���F_Jf,
&�,����t�􁹔���x��I�~��L��\ �v	K���[�2^����,ڻ:���u���UTB2�(�JSW:��ȱ,�����{0B�L�<���1��Q���-߸+�\LQ���q��ÏP���`YC�e2���8�2I���|�a+B'��f�Z,'�R.S�V=��`d^Bqx]W�@�M~�"�z�ozY&u����=�nYP_�	�n����6JǒT__'Ǝ��5~���1���'�{�yx6�e8꠮=:�a����t*+������2�X܋�c�b��b��([�O��*yP��K9nv_Q��j��^�m�zj�0��?�X:��ә��Tt�=�8=0�Az�WhԨQ~��\�b����
�w��5%����C���x%<�x�Ǳ�ι��m�����ի[i͚54w�\Z�p!͟�6u'�yQd$��yi1"Ns��n�7(W����9�h:��i��0;:���rCǨ��EF�=����V�E2h ��jذa��C�]w�!�yZ��<���	<�ޒ'�)�q���.cuPl{V2�l�Ϳ�?�x_CALD<�L&[xcySʹ3h�IV{�1��<
�8hD�M�I�U=��*�䋽�T�}x&�L�I�"���_�/�.��j(M?_�g�1���矧T��
Ā̉���]��X��&L��u]y仰Cϕ�X�k��T;�&5g�1�IS��u'�(�|z��y��k�ѳ�?G�^z�s�M������#Q*&�<�������r1�wwuSmM��nt�q'�u�p��=[^��,��n�/�n�Z���z�_x�ǝ��H����׏~?~T�����l�;>���Af�)n��!��.s��ˋ����#F��{�B�I�Z���2�w��T��S"00�i�XuR{g;'���g�^J���^���keщP�P0���U"��^��Tl�F��sS}#�4m:��޴A,�<� �s߽�}�ч��e%M�4�� ;�sD��*�^H)�����󬋑X��n�{�ځ�sa9�Vu��/��:�q}�����/��<9G9'c�no��Lr�ر2�.%��$3,��z�z�7SKC^dW��Ȱn��g_��~�<X�e�ĘFȧ���(!e,�b�E�L_+�B�������a�5t����	�q���]w�Es�̡�+ZأAn�� �cZ���֪D�}�d��[藤����&ߩ�����s�q�S�۾2�՘Яe���q������_���I>�����e
-27��F]����K,X��N7�knC߿�{��N;QZ�ۈ�3D��j2�-��y}d�;���@H-V"L�a-"=/�KқӒ���_�2��^�����~�i�-q+\c�*Y�Ê��c��b@���Ɏ�V0V@��qfWf(Y�`�?�"�r��;*/�M����d�5ʚ~K&0�=��>�#-^������E4`Ճ).�K̘��oA{:��׀X�0�mcc#}������1f[�R�B��=���g'�7��a����]/�7��R�����`�ǔ��v�CJ�}�ߵu�Qƙ-��$��E��yԖ���E�N<O�v[����F?��O��o��m4z�hF�Ec5��Ŕʙ�]fqD�<`8~�cO��_�k<k>2����pM���G����^6r�%̃U�v�o���vT�2��ݴ���R5�Eƃ�s��v�6-�
I���S��"���
x��.:C}�tgL�����/G�&t�|��U�0"�B��0 k����T��+X�O:�$:�S�o����'�u*���L���6��.��;XqL,�@9%���P@�566Ф)S�y\35�7Pӈ&~��ae�X,�b�F���6����.���q�/iժU��ȉƇT^��P2����X*�p��s<^��@�,%��3NLCۃ߃�[�l���JP�$9C2��)
����pۖrŴxHr��hel@M��K�r���^��j��-1���gx	��~�K_���;�+ޖ��W1���,�}�l�8�W��w�}���կhɢwȊDك��J�7U�'@� ���A�;��D;�Yx!�h�d�pƎ�[�~{�M����ے�s�9���q�|�u������ӟ�ru���xM]�R S
�r�*���s(Z�Q�FR�8ư�0�c?/U��0���S���d>�e��h�w��H�4#���q=;��t���c��K%1	�7m�e�$����y��=��_D�#�1����ӢK��A�ȑ#���F3�����Jp.�r��6lU�P�]�tc:<�_��Rԫ|b�t��7Ϥ�c�p���P�K���$��%< "�K��{B����	Pl�@��keHkŊ���8,�<�oS�H�y�]�k'�@�{,5���߅�q��u���MS]�g�}���::)��3�ַ�܏��Gc*�qBY��������_*%��a�l{.-�d8��C�RJj����/ж�nˠ���$?��Gp���*�={6��^C��O�*��ČN��.�EK��%�� n@��)o���;�.�l�E����̡9.<��(��&Ӌ��Ĝ�%.������ I�dGC��U�s)VkJ9�Z��E���V�9���������@�:�]�3)�#� Ixb��� r�"�྇y� ��B(&*,�-�#'Il�xT<y韧�-� �xFxAx~i�\Z�x1=���t�wΧ�g�6@���^3c�(��f�����3Π�-+���^��	㨭�#�{�xJ���z���0Tc1A����b�?Xj�Y��ɀU���tnNsљ�}ݠ`#@��!��N��f:;�+B1_��Kh�i;�sQ�I��9����g���q�]�~]�!�Hи�6o���X�M(-q���+�.PT�eXַ��ji�l�$��q�<�lzɣ���V��-���/'cs���>*u���7�ɤ��dW�ߍD4�c����.)�ݓ�>ZX�G�&�~�Bg*A5bъ[1�Y���}��� &�+�>���	Er,���_��Ï袋.���:*�8�(�s�玠|��[���V��{\9b*M�����A��A���%�d"qU�j�����f*M��n��4cO:���}��<�ԋ��i�������/��{5�"���'��Z��{�1.�&$Ԣ��̨�a>�B��2nu�l�($�º��h��;�~���dshvvu	k�����������Q�F�����I�5$���4�F	3X��c����~�^~�e���yۯE���5�;��;�����oм饗_��b�d
d������wA�z('W�x�����r&o���q���-�K"�%�Cm���ӟ������m�r��⫯�F_�CZ��LIRSWKV$�R�J�H�\{���/�����UV�|)��7���a���������l⨄+�(���v�}���^ȋ2��wߟ��T�~��y21�[,��?@����~q.���=�AP8�X��f��W��Q#��A�
�+��{�;r�!4�?���Qԍ
���$�^���D��t���n�@ر5,RDx|0H�֯e����z:�3�C��\W��sR���}����wߡ��Z8o5�ڂj�k1��c�*��ׯ�W �f.��@���k�,O�R�g�W+���I����ˊP7X1��`��8��C��R�<sl/Ϗj��`̾Z�50b�쥂7�y��"��G?���t��KX���z��W�뮣.�.m-�Ir4D-^���U\=走��b��Kz��$u��;��blޟY\�!��1��R���;q��װ�6o�|���WӬ������	%E�0"�?�����?��:�vF��ʥ�<�Ś��e�N�x�z"����I�\L��|�l��� C�5�׿~����P�^p��aܐ�*d����ʫ��_�����VnQ����`�Z��{���WT>ƺF�!|��<�F��� ���ֽht�7��D�1���J��g'cU���0���8;;:i͚�4q�	t�%?�O}�S4,���0HjbH�&�K/�ŋS����XSˋj��r(Z
������~7*L( �xQ}��'i�m�щ'�����F�"Ž�ދ�>�h��i����d����\��0T/N�wa]qi�}����;���8��o�
o�)��믿��~�,>����ؑ,}|U���A��b|����:��4f�X�v��d���ՠӂ��e�(����3�;)�2���G�T1���++���	��T�D�ƌނ��ʱt�	'�Ȳ��.�uwPmM]qŕ��}�i��1F�.����+B!Ϭ��;깘�����n�\��,�&��CX�P�`���n�:������N�5ӡ2,��y���뮹֯�q��(��11�L_KV�&����%]4u�����8��n�D�[WR��ZY�ʁ�!=���t�_��a���)	VR���(В�*�,�P�bz�P.@�"d�\<�S�7L�j+���Y�?}:�������Lzܸq<����Mm\��@�v�2*+'�КL���E����Cx)q:����\a�FB
����w�AW_s��(ӧ��qm���u�AU*�T��I��=^*�Vs�`q�������K�?/ͥ�!k,�g ֤(�'��MM���d��Jg� ��X�|������?��t����ƹy�5S�N��晌$�����p�ת��A��H�9�1$������L��cƌ�:(�d�i�M+o�7�~���G��;��뺹*&���=e|,m�0�QFAU��@��㜇He�?LǺ�����/��&�C��j���y�./EO�y����k����qf�B}Hcc�o�C�"��G��C�xߓ��SH��R�r�g�Bu" G��H�k��7(i^x�:B(�Na�Gjd��>��D��M�F�~�3i^�f5���2D��Nm�[л���F`�'!�,6MÚ��Qg[;}�����?�jmV��g}{�l^����Ut���T_��S�s����l��Q��i���6�%�O���03�s$7�m�8��<����nX܀;��P��)���#Eq��W\)]���%}]����BC��͘���w�����T}<9� ձ1���׾��Z[WѤ����?����jk	�\C�P0���UWq�.��TaVn'��]זw��Y%�k�QƖV(���`>M�qZ��0Κ㍴�>��Cb�����i��#G�9����O�J�}��T����S����R������[��Q��2/P�a61QP2|x�3\�9�hBgZ����"k����?d>�
]|���o�y��CU\�b�N�I�'L�3��M:�HYd���w	'�Dɱ"������y�ihMM#h��u�:>��D2C�����
H+"�|tĴ�M�b%#����z�A��}�%Z�d1�J�[}��t��Fq=�0n'�7t�Iv[���*�����ĕ�ĽG��g>s(}����|Ӝ�xQ}���&R��pc;�%ʩ�������-+�D��b���22Lvw����m���7W��yo��teіjjS$S!2�*�+�P;��Iw=]���?��1����}��$�{�$St�-�Y���{v���:Z�z5��`;�#��eS�B*�Dbi����P��w�4Ec�f`Eؘ�;?mmmjA���q�t��gSC$N]n��v<�=�Ҭ���,���Z$S��،k�)ÛT��g:t�M�r=-�ɓ'SC]=SF ^�F)&T?�2�ǓJ�N�%��ci1#X��`4= �CG�Q��Z �����h�R�gw�,�0t�Yd�~!�]��rAU*E���?�.��R�ޣ+�b�X���k;t߃����L�W,�ѣFK@�XXŵ�,�7��Z�Z����.p�ŏd����U�^#µU���=��2�?�s��.p}��?7k�H�Aٜ��~���4#x��ds8̗��.��Î2<Y@�q�6� G�l��2�Ef���V��o}�&����&"�yvIq� ����9A�G���������~I-��N��^HC��5���E����SO<��d_3��l��W>�v�.�uS~1����~# q}���ٰv�|��ÛewH2!Y���5��v���^P`��rM+�Zf0b�~3#UA��g��U훫2�~*�40/�43f��ė��7��AX�	��� D&��{���o�U�x�R�Đ0�LxJ&1�	Q��Ғ�.G(�d:E�֮�D>�o��IHwF� ��d��+����sy�'��q�O1G�|5�l q����v��ꫯRm]-�O.���<��Q��V:nF6"T�Ϡ��"M4S0������NS�ߞƎ#?���4]��������;�̌�---�j˼Ve62�A3{��0U)e��t��P6&L�o�s�>m��?KL,�X�K��f��7ߢ���%�I����aȢ=۪���L
���
F7���Ba�ʕ+�x�P\�@�h�xT"r�JIo�K��-w��'�5A�l�+�a\���t�]w�{8o<2�of�S��d�?�S��
�ٷ��G헛��Q�4���JG�ٳ	Z�ny�Q��n���8#J��_��f�
��.S�L+Of�ҥ����E�'p�zZ%��b�E"p��I|7�����s�	�9�Lr���SO��y���ύ19֧�t�7��Y�h�ĉl��cqJ�fɼM�C�g�P��M���U�$iX�r��B?'$��v�؛�F��I�����&
��-�w�+C��[n�R)z.��*��ӧ��_�
u��â],Zqq��k/�?_(�aT[��a2(cx3N Q_uu�JP|Wf�2�ȞI��3�*L���.$p҈j%���4o1Fޥ�3S�����e��~c�����;�8���^�=Γ��'bd}y���E�2c���@s[�\��ZT�wז�Ll�a��As�����/�������Н���?���{�&�z�1��2�N� �pSث�(����͝�h�B�/��g�38�J��|2IK�y�~Lh���mY�L�����/��ѿ�����ǔJc�>s@��P�|��E�kl`
�{̠C�4��A"���k��3�>����#�������3
a�}u|��T4C5�2%�(s�i�}�t!�nJ����U���f�� ��L�a��[�[&wty�j*�p�9���x����T��1s3��@nՓ�?q%��L*%,��v��sG�9�|�j+@4�;P[����,�z럩eEoj��ߕ�È�$<`���ȼ���v|߱6�J��h�N��L��o��J+�b|!K[���"�zi�P&�irrXX�5��k�Zf�>���;��p�����B��1��;�Z���'�,����@�KP�J��CD(ɞ���ȏ\	E��\�G���K����aW�-Ît��gfg-_�+������9�]{�_d6aĈR0�d�ȞH�}�4�qۭ8�k��d���?��fN�x<&��x�P*���gXL�����8�:�?�զ�`Ֆ������H��Y�h�me?����ym�6�ҕ�E`g6ce��_�m���c����c@���ɓ� �9j��a��N�K��ѻ���u���N�qI�Os#���O��`6UO����m��^�=�i�s��U֖�n9L�N�x _��I��ͨ��E^%�=Ĕ�v"��)$����p��gq�b�e���(��PM�k���r*r��ԝ���j�A���_��^�MN��E�CW-~hN�!!1�آx�Pb��qrF(�]Dy0��>/7��?@9un%��͝c������ŝa���H�:(a6�^��=�g�q$-{&�0�e�?|���bp�� x����4G
������������0��<��_5�;	(n���4b�����6��w��m�-my�a@���` fſ/'Nd4ɚ5k|M���^�jìc�������`r��'����>����B֝q1
)�����%������P�y�T\�kB(���v�����g|�t;$�p�ס.F�/x0����x��Ce��x�eYY�I�#R�â�H�~	G6!F$z�o2`���[��� ��	m����se��^�$����15c1^�����q*jF�bC�:��27Z[9���+/β��'{�'�=>�n�t�B� ZW��G�P^�@�iS�]Br2�h���Q��<5!(x�8o��_]����~λ (�^#�#(������T�l�K��hoa��LP���9A&+�d����y� i8�ڰUԬ3Ѷ~G6v���U�I�?G?
�%��<?A�)��3m����pLd x'��� �ٍ>I�
5/+%���~X�lnb��bAK�����Ldy�I'1/Y>i�G���y�Xm/~�B�3�%�)����U<'T78RnFz@iX['���V��.�\����9��ihl�����(�	�FG����#�Y�.��;Y���?g���͜P�l��}�����v)%�^g<������7��~1?�4�ʜ}z��~ƌk�����j
�t�����;�@����FR�c�1���u�s�:0�<����i���;z<BIuttp�)*i��J^%#���/���`t/>J��5.�ފ9��#v� ����G����R�h�
����[(�B��t饗2<9b��G��8s&�X��jG�$7"�ičp m������I�Ն��_=���~ĢIr�8�Ϣ3z��m�%�M�<N��0�7P�1��Ű�QM#�~7�9dղb�O���E�����6��;�D\p>M=�$��
E���a?1���¾kԷ}�):����@9�*�SU�o�BVM 	��"� Q@�dDa\XD��:��8 "�"茨�Nt@e�EE� YI��Z���{N���~[���[�`�y����Uu�w�9����g@�5�h&��2{���>@��'��2�p^{��h���D�P�|�a�ַ�e<���y����\R���5T�#�*�iX�ۯS��Y��W�x3{��Z�$��/]���Z�m�OxR2̹��Ƥ?���!�¶�l�� �¹�-�O|�����;к�njok���|U��_�����O}���.$�A�mV�e�d�A�NLU0������s3��5��hYì6����2��
�d���i�r��˨r�l`�!!�U�a�u�\��< 4�ۚ7M��?�s�֜�(�,Km���� L�
�n�&%rN�$U��jc�
��B�z�4�m*�6Fh�*�8�L�9Tm�,-�'ק�\�8�k`t�^����
�3@�Q�ZU	�ߺ�¶��l1 �Amق���ɋ��yݖ���+4
͵�s��BO�k����t�s��W��aIn�Q�`��N�_NB���k����Q<|��k��ܪ�����9�Cx wlD����2�'�����W|��2@�2{�]�8@���@����" hnzPh�$0�^(�
�u9�f�J��m��q����ӱ���{�>�������ϙ�W~e���[�lV��՜����a�e�ٽ�S[���͛��(�� /6�sWnfM����+y�$�a=V{|Nz��A~�:(��m-L1���a/��7xo\�טڬ �����Ё��O(&�>��g��������H'��a$m�y:C���B��i.k��W�D��~^�D��!'�BȄEe����gW���s��C�k��FFv�|P��d��x�w����u���̲������L4^��m`|�T��%+�U$V�H�x�+��w��'�M=f%k^s�3�N���8��.]ʀ���[:�5�$@��͑��)��5tǃ�*h����t�}X���>�Z�b�� 	��d�?��G��'?ɱ���V�vƃi��y������\D�jl ��l�?�1���w�e�n�,�N��赵�}�0�9w򿅽�u�x���t�GҔ�)�pZ2����V�n�D:���Mͽ�)=��nx��S��ş������^�2<i��!�5H�ܲ�-^��WM��w���M��3��UP����.Zqb���r2�m��L8akV��� `��m<�2'�a`.��c^��>��Tϡa{�5��@���������#aǺ`3�,~0IT�K��g͚� ��ʚ5kh�����ƞ���D�u^`J���3��x$�ꃹǽ�x0?������^?4|�u�����m�Rf���*�����w���
�����7Q+��|�3�<�(=c����#�~��������Z��w�HimI�8��$K����+�	���w��~��f����Ν;��k�M���o���.�9���}������u@S��	^�77�[��^ �y ,𲉨Հ˦�=�ۛP��f��[�%〺k>��S��;� ceު�ו�A�M�m���{�-��ׄ	�m&qs2~bWy�j���f������R{�sgw��x2h]�^"�jU��۷�OO�^!�dx[����}�.��픕=�����������ᴴ|��d[��pm��PO���.Y���T"7�x�������Xaˠ/����J#��̓a�!e�9Hj)̖fK"�s�����'��F�Ӷ�D=KH���vx�a5%`2�H_�Db�j�&��8�0I������0�:�����]���&�k�D���DkVo��6s,q-�@�_�������J�˴�Ǉ�T�UC�n��EL��v�*�ՇFw{1��������K���?�r32=,�n�ì9s��D�H� pӼTl�?�ir;��+�oƱB�a��f�c�{'���no�Ș�б����b9E%I���rS�L��?�ܔа����|O���������Ti��j˗���tcr��;^5���o��=��sY3e���ͼŒ���ib��L+N©��X^��@����7n�`��9��c��\��ӒE�8����i�C����qh�Z&OHj�V3!��}?o�Jgx��	�fv���O%�1��"
0nΛ��W��m�c*A���O��L߆�z���M����rM�c�E�Иb����O�S����F\��ͣ3�8�v�a�zi�*�1x~�aN�#�����Y�q��kGd쎒tq�Zdl�c�=�@�X�z5͙��|W?��I���B��/��Et�A�����\��w��kn�=�  �j@���i<���d5�i� ��AA���wۍX��*�����i�}�Ӝ9s6��~ӟz�)G��q�.��8�&�maf�2��ZHǨ�z�$� ���T�,bOEV�`�'>{��<���t��	MyY����0��B�[kks�  �)�%r:�L�5&S�;hӬ�ƫj��ѝk±�� >�c
�]���\���?�xu�j�����?�}�s����D<U�� �F���J�pC3��D�&��B��<;74Ϩ�xD�N ���dԸ�\���؝=�PvF"���2I=�~=���>���^�:}:6zV����!��76{��#\Dm�=�/�����enP�lY��7i�v�f_ ��`�e.����������|y^�ka��[���ċ�-n��A�f���v�߅�0/��e���T13�ӫ��?����}��:�+�� �$�Wc�ǣ��0*�^��ל���N;����g�?�z�'"ܤ #��$��N�~s��iݺ����v�:��|�1%�)š˲؉,��FM3�ڿA�^���4m����s���<�"��J��=d�������"T�}��]��f��6Ή97Yè���2�L
�֓�ڠز����X��em��r<qkn^Ti��v�4�Z�BX�d���W�b�j)���>*l�U]�m��|���8X���B��Ƴ��l�x��r�)��K��f��RpI�7�����0�m�~!���dr���.	7M�1�~����#�?V[�Y�h5�{�u��h��uRR�����7��͔˘�Z/l�H���O����ٳx�SYz��"�9�ujz�z��X��$ޚ~�ꅥ�Ps91T�I�a���̦իiދ^D��lZ�x1��i`R%��3w�w��_ߦ)ӧq��A>�����ʶ�2��$�U��}U��:��¡��V�Ǚ�XW߯4=���&�`�*��y��[F!$�A�"�������?��j7@�Dp�4���-g:T���$Y��.���;���Q�z;������O�gL�g�YErl5�h����!]�Af�]w��$p�A���u�c�ꮮ���g�`R���E\���3��ݰ.�`�^�gռ�d	o��p���EX#LT�Z�A�LT����q���B(�\=�}�v�zz��'���%���*G8�3-e������޷}6.s,}_�9,�UY�m!;-6�w�-�7�_O�����+�s�t���qB\M�W]=�<.�Kn��v���{m8qJ;'�7��,�n5�`Ƒ�b�a���>���;`��.O(�5�?{�1��dy�R��g�N��{R�Y�b�8���t�]��֭^G/=az�g^?�_D�l�*��{%}5'����(� ��#�9Ȩ5��h[^~_�sr3��J��9��z㘿��Ą���Fm��4t��/���2�'B\�,�p(@���iI鷚k��t"m�ln��v�o���T���YIc<>n��V蒄�=op93���*U�*v���z�\!����\g�Ǿ/�S��v�@��w��I`"��Y������8i3^<>O@������u�ߵ23�I��r����c nڼ���9�F���3ϯ�Jn���C֭����t��6��^��0���c6џ�b���`��;��<u�N�ͧ��/X2�۠@�����<�l�ǡa��%�X�;���p����L��+� ROFz����a��w,�)�d 2�u�]�����|�5k��G�De�O@*�\�����L,�-�T��q&J(��(����k�e�VB���3�Z�>Vt87��gӑGE�>�,z�+f��� ���0����ѣf�_2��b���N�%����?'7�����՞5kh��w�]_�k�����-���~���?ta3N�&�َ����s�3x.�U���>3z���,�v~�N\��:*=��Jt�	]���2��z*�������3fH3���@��3�C���?�O��)ȳ��\⭢y4�
���Ÿgw�&��5��Bu�_���S��> 	.r��!U���nI}����w��W�*x�i��^�On���\�<j,�h!�lfN�^>���\
.��#t�zz�i����h�Et�?G{�7��>8 o �z08� �
���Qn�˖/�0�!2��e�i֦��������D���u����Rٟ�����Ν��$T5��>�^^��)�k�����u�7��uǓ{�`�Δ���0�.R��6\�8���������|wr��Ouׯ_Go8�h�>6�L/�R|2�n������N�~fP ��.��/��6l��� ��f17}J��W4��Ab�9`��3����t���l�%�*h?�9��������O�d<��]e�	�'��˲p����d.\��n�@2����
��3 �i<���fz�?@���ߡn�wG{Gڲ|���0�鿷���M��3g��> ���)J,�����F�4<����5�A�,�����Q�[MxL���/iN�P4��nP ���H�Z:����37cB�z3�@�b�?<v�|qݨ�m˯��~9�`B���`�n��O�S,�`oZ��W��S*�}�ݬ���SN��
��0H�z���S
��K�
�ܢ"a�L�M�F��������ś�d��n3Iϲ��9�*8�θ�9���[�	��o��͟��2��g̟��g;Yy�!�j��/ph�,��iܫ�6
p�׭ ��D��vzա�һv�
%Cϰ��L�A0�s�?G�<�q��3w�R%��mˌ6�[�Mㅱ���MayS���|�oo[�=�,|*�,rh�9g�c-J3�U����LJ�E�ϬYMW�����o�¯��hs��2�H�v��oK{F͜1�=���ſ��o��i?r���!Z�����ҵ<�J�D������X� �ήNAË�>}:�>��x+���o��dJ'�p�}����_��̞{�)?̷�|iˌ���Q^�9`]�l����H�@^K2��{1��m����ʨ���^8̲|�$��,��In�G���v���������[y�V&i[`V�U�v�>P�n3���m~{��t�UW��߹��]/b�2%���t�|rR�)7>����`����^az��]��8���n��K-�=aT�]>�ߍ\L�nm�"LNG_6��E�&�|�d7��FzB[&��\�z�1	�y"�`�:�l>����^D]�7��X9�y�w������`����re��{E��̝;��s�9��7ތ�5nL+-3pn��i�*�(�����2�õ�L(��mKMYnzת
2�kO�/7�!U�������_�������Js���N�iQ2��p�3�[�(݇� J�Z�g�C�%ͳRa[�jddr�e��ؚ��6��>�S&�x��_�	2��g�ʂ�=��1h�w�s�Cф�*3�d`�p̀���w��
���>���Y\Q %>��x��N��i�z�ys��h@>��ߤ[}p���U�I�j�¹�M�]�����~I�����_��W��ߟ���c�,���ޞ��Q��Vۋ$aԽ�F�T4Vs�M;o��skV��"	�YO�H���)u9ki_�����<I�Θ9p�Z�1�a@R��O�.D��Y�p�S���s��ɮ�j�҇`C�{ｹcBf88�ii����-�7�"��T?��F��T��-eX��A�VE�A��]۪���)74׻�.��L@���e@巿�==�j׆����w�M��򦴳 e[�����SY��j�6nsH��~C�C����ɨ��x&I1��E��	E���D���`�p�Ϭ3^�K���0�L��uК�kX��uG��~���z{��ܖ����VZp�3 �2��w�W$?�����̙3�������o���y�(���,�;W.��*��� ���Oss3.и��\����M+)��5��}��zs~�Z��9_��1�L���[�%{��WQ`���_��֮]��N�7e�'=����õl*�P�u�]w���~�̀�nS�W�Ū�0B~?�3��i�Ř��Y�z=�{a=��!�r��/��!"�͂r3M�a/��Js��W'��!�>��}��<����w���F���O*�A����?�U�]G��x�J݌Z�Y��w��������=Z��-b�M��p�p���TFƵT��ar�-�"j,�P��D�ó�>0G�ŗ�̻�zy,�~��ft^��vfW�S]0��92�Ky�z��ي~ϠAf%�������o�|��x�� ^Ÿl>�t&�no���7V߆,��p���D|�g�K�ק7�x H�x�V���U~�b+�ďX��?�)��'?I5z?�c�\��h���RX��3�PUG�)"jY��p)�o2BE�m�m���6��]k6��@��`�����i[���ζc�Ҕ�/�)I��S,*�}b�=?��5o����㸵�����e��N�x��,�����8�X��ƃn�׼�5��C�D�A���Y&��M��Q�,q+k�5U(dfƜ����m�mY�=1F>���9�U�j�\�5eU�}Q���h�j�y1k�[Eaǣ��7~��VOM��5(¿���ή"}${J��=�j������D�3ꪡ�^����Z�6��� `��PP/l�*F�7p�g�*��?�ޟ�j���9ԍ}ԦW�Ϲ�ϥc�y#��?
�6��,��>�Al.Y�p�w���']t��G\�2#X}r���/7��LJc,?=1:a4�����kLw4�֎f�6����,��T�Ia$�#[�?K��y|,^����eWcvU�X���i����A�W|^�*���Rt�:Ms'#�y�s>��(]8h�B*Vbț0�����jZ-룏y�ĺ{�kd��*��|�eQ���>��CK�.�o�����`m( ����;�Cd�f�b��tS���yh��ff�����Qm��o1I������v͕�h��1�UL=��#	�#<�6�)��?��P��\�!4�2��q��6��O�DZ���R��$�ٟ����y���rkL�ޚ��z����?�F���9T��D�W���l뚻�ST�0�T(3�2�L\_�O�$-l��y�-93�r3��ּ�e/�j����V��zhm���!D�4T���vV6�ꘉ3�8wl�Z��ƚ1/?���;��-�����mhq�\"۶��Z���4l�nZ'����
Ŕ�R2�KBV���%/�W�� ���w���{8�4����;���t�M������M4�-˕�GJ^ pK<�%� �e1�LZ�V�&�~|�7��J���/��s�<�cLY��	涶��,c���������BڒeHvu���+_�J:��#m��[ڠ��ox}�ӟfo���-}�akd���gTU'"~��HBn1�&3P͇+
���6br�c�6��NJ&�3����JH�74tFv�D�r�%iy�o�lB�v(��n�v4�%�[
2=����^��W'O=�wA$)���srI0E㈥7�c'Ǘ����G$��] M ��i�&������ms㾰|��|�_�lج��k��Hp��ޣ�FBg,�@�m����j�}��:F��<֤�?��x�܆yј�>G���/ߛ<����P>�5��~2}�{����i�M��B��N����	�y��V�x�*����o�Z��d1WF��=y.<��&���
K�@\B�#�_����c欙��giÆu\|����7���w�mf�]bw?R�gX s�[O�9����K�f�fZ\3�q)���G����WA�Xd���s��}Y�L.+�wa�\Y,u[u �$u�s-S��E��e ���˶��x3e��, �4w�\Z�d	Bei��0����������M9蠃��Ga���N�U�R)���;g�yŤRXa�M.�;7�4�EBc���q��ԃ ��������!�#�|-�����֋��������e�'�=�y����7��-X��u��ո�=�$��@�,���{��Q��7���W�4Xb-��o �F��+l,]�Ç��֬��ㅍw��pÏ������ܹ��eZ�Te�����Dt�<�O�2�K{�����ih��U��;̣���v��sJr(�<TY�-%������,/:g��?�	+�"7�n�v#`���8p�Ĳ�#ʵ h$�PXa�6�-�ei����3t��wLh�ǐ(m�{1
0^
:�������n�}��'x˖Q��^��mɒ��:��Q�2?l���s�?���˴��PwwW��+�W{5a��[���֓	q� �ӎm­�α�
]���\�B����b��mo�<�L��x��.�@��)ʢ��z���/هϱ���6��
k���t�i����C
0[ӆ��'	.��eS.8�M���-4{�,.�D��l Ü���!�}ȖT�^z�`i�QN����
+l��z2��:e�)� a���d�Tq�Qb��V��|yo� ��}��s�?~7�d8�5ߖ�L��$����_�|}�s����g�a-$�'��ʹR�駚ey������7��B��D�-H '��M���S���b+{C=���o��x�=�m���5����]���/�0a���"I0��U��IWS�=��p(h�r
�V�X}{��7@Y{ݺuܪ�㎧���ej�W1ӯu0�R'�ڒ�[?�p:����G��^3͔���LGf��h`���q?Vu�<���La�6��Q5�d��j�Kl�e�H���1���2�dHe���/���>ڀ���e�x���Th+ږ�L-������t|�O/�Xג%'D-S{{�$�Bd�P�!�V����(� c���J9N&�'R�ĵ<��5m�Qc��%�[fYփ�s<�Iq�b�;;�q��*���	j��'���x%��j����d`�W�Gq�w�!'=�0{3mm�2��\��z��v�� �n��c$��-ʄT���AN�8ih�J
+��¶��Cd�Ի��8
�
-S!bIV�s0YC?��!�]n.���>J;�#|��$�L߅½��d�ҕc.'���U����^Z��t������}.=��������B�J��p����6���q���Ii~Fc��C2�s�U{��Ma�6V-�{�DN¤!2�T�L�`"4�8l2N���0�y53\7����	_D�����c��ʜ7^�"U]�"��d�k$<��,*�mV�Q�o\���������.[ T*��e�Ğt����Y�J+puP��I����Y���
+���d�z�T�1�� k� ��y��_0Ϣ&���^�qK�wܑ��w�������ߡf'�؆MaF��Jz��4)м�k骫�bof��M���5s)���XZ-'�*+;=������_/�-r����n��앭m����u-)ֈuV*q�����Js��NE�P�dl[r���&a���r��Kk׮�w��]t衇Z��Q��L�	��Ȃ̙g�����7�����;�nz9�5�f<�^�M�^ʪ��'ߞPKe����W�f
+��qf*!I�>��Ծf�O�m�H
8� w��h|��U�U�T*4e���׍7ވ��p���|�\�ђ�� �@t���!z�W�G}�J���;ٛ�9{��O�܌z3Pm������oOE�Ƿa2J]̐�� 
$��fKm�+��N��|e?�a�c��&�����4\ň:-�$�/�����k�Mde��\��jT�I�Ӂ��7D�/�m�S)���;::Xm������7*�0��ȁ �[j����_��[��~�[^�
����\��A�_���O�]���y![����dO:Nf�Y�L����;SXa�����3vƋE���0��}?�)�?����b��3/e�uuuq.f�t��7��M�K�,Ќ���(��~^@��n�+.<�����ҦM�i���}Ǜ�m�+�wZ�sޜ��҇�����C��2M���|�>�O��d���m]s��9S  �IDAT�Fj(��o��oiXL�*�Ж)I�8��wɷ��̮��b;���oJF��>� ��YL�KR�(K��ȸ��ݚ�g�qO��K�T��7�Nհ��7cs3ޠ\T�h�8�Ϥ�1�R�u~Na��ul�s �H+�ON��JǸ�~�����P���k~"@�|0РF�ǟ���ۗ�?�|���ou�-G��ά|�W;i�W��i}�M�[n�&m\��usZZZ�7�5 �Glw����qM'7�&���s�Ѽl�h��9�C�!�����_x*�mE��K=��v�t�y�L�D�R`�\��H$��̑�sNxq�?��fC�Z0�yv
-y>?�f��S���;�������JY�A�G�Fd��Ʊn��|�=���p�'F���M��okk���~�U���f<���h�I{_���C]�* �LP�f
+��1dy�#mg�UVVN��F�TF&�H<?{LIU`�|���8L�֓�J����h)�,Ƞa̲e%���2��n8�J7�闿�%�Z�M�>�Oww�-ؔ��ǉ�0��x�
4�ERH��(#�����߬(�k}_��
+���0�阂	��jU:[����g``�T�����7�Y�̝M��-b�c�2p%t�	'Ы^u�w�4�f��M&���|�l�򘖓m&s�}i�=_�}�K�/�f�9s����l��dMvK�J m�L$��ښ N���g���
+��0`bi��o��	m��qѥU�ʥb��.S�\�}`Ps�QG@>@��7߼�[S�r06� �y�_�>���w��?N==��Ĕ	5C�� 4�y�R�-�[��H\_��r�M�����gFFĹ ��:h��< PC��-���̡�7��Cپ��e[����y����}�6h|�5#|��`r�I�$�l?{-BQ&��A%�x<���z>�e) M&��s��l�O6}�L���]�ژw��l:s�w�\��h�y1�ѡc���ms���]u��	�N����e��3�� �ت P��+F���j��}Bp��H0$TțVXac��y)v�'�>Y�ԿY`{x����e�z�W��`�z@e?:^`�;�8x0�(���ml�2߽?4���KZ�y��������	.75�܌6��#V����^
X�&4�	 �{��%�e,r2�V�hZJV�3�2Bf�@vD21_��T�Q'0����r��UbѾ~�z����?H��~�F�rY�mmc�A��6��?�������z�����d�$S�8{�K6��b�ި��VXa��
�y��t�Z$r1Jh�i�?���%����������Mo�f�|l�{0j�W��~3�����7�W_}u|�WRd�<�o�7�r3@�HNn�ĀD�s������JA��q��}�j�֊�Ka[�����h�������$��Ἃ�U�L�?''S�?O�,y�4#=2�R�v�fΦ�}��X������[n��[>=fF�h�����^G?��Ϲ[ܼ֎v����f�'?�I*���+��LԚs���
+���0ͽ��M�kc� L�*.s�:�}�^6C��(�DDh�w��N;�n���Q�%�m�E�y��~{r�y�@���|nF��}�E� `X@Ss:�p*�|�qa�V��2`��J�j �b7� �	�~!��T}�e��`ss�m�b@�H�u��~G������m�&�۶��z�q�5�������w���n�՛I���0�(���w-q��p�&R��P��i#4���P)ą6���h�V+���0������JR�#�yXF���L�E���=�i��gδ��Jwϛ'��fz��|㭴$XN��z�cȶ��$T�:�,�뮻��g��iӦq����к9)�)�B_�^k:�a�M���-��&��{17I�ԝ�4y,�� �y��`�Os�}��u[�g�~0}��k���eZc� �+�d[6�_�6�"&����o�6R���������N�a	 ���O?HcͶ�0	�/}����~6��?>GO?�M�>�6m��� NjE�K�-%��VGN�8��8(.�/9�L=�W��%�� - u�`��V��.<���:���&���3O��r�s��
&e�nKJ`��\��1����������o?z�;�A�\~Q�y4�ߘ�?�V S��-�:�[�W����~�?\��f 	d��'�@�0�{�s�,���p^�P  ���5ڙ�M C�\����ku=�11�Lxk0Xs�?���bA؝ӈ�.��Y!L)��^�-ͼ����}����h���ö-@tl�5ϥ�;�������;��̘ �����%��a�ԇC_Ҵ�1���y�3�$#_�z4�E���[�yN��¶�Mf���]�>�`�+b�z�C>�c³�ecr�̉��T��,?2͘�7c-�`�*��f�"�]3���/�{�{ݕ^ڼq#�{������m�<fm�x2X��T��t�S��tӗ�g����6fc����ʺ �CŇ��z��T��Y�Xh 4�@@�=����S/dnCZg8�"�zqx���*��բ���Xc!&�^����a�#ÿ]�ɷ O�H����4���<F[|'��/jr�w�׶�s�~��	��o��{�<��I;e�a��u�J��E����߇�rX�Ў;�D_|��[�칍̇��D�ll����F-Y�|�k_��կ|�vj݉=����J��h%�+�P�jV@N'��Ղ�l���(ų/j���$���Z��4K��P�oy}�\7��%q�&T֗��$r>gp�& �T�i�`�J�մ���qے����H�%���1��L#�QϽ�ג[��������W�2��/_N�_��K��4�m[�L�|ۃ����Mz衇诏?NS�Nej3Nz���7AR�Z�g������k��^F@x`�v��9�Yݠ�
�k6Y�p�*�@������e^',�x@ 0GW�/����,�-0^ �ʳJ���2���g�񿱌rοҗq��o���>��'л~xc�?W�#����)�r�Ɔ'�Fg+V�/�{�ƛ��\z�Gxe��ks3�dc�����SK���O��N�&��R&-���Z��\�����E &(�����	�h��]E'��(�6��sў�g� ���V�b*���c�H�T�߿���-(�{�C�Qi���l��΢Ay�����Vk�_M�~�bz��O_�k�n(�����ZI+���l�d��B2 ���:�t���~w�r�J���Z����rmeP��1q�'s_�(nb"�Ϲ�2m ��2�82�f/��y���.��w�/�:���|�$��,
�f@3q��}>����7�3��ܖ��t�CY�q��f[�m<�r��GB6�W�ZO��}�5Q=!�@B/0�J����AL�õmM$����h��-�Ũ�B��������޽�G�d��h^ͧ3f҆��ڴ������w�;Gz˿�D/��ǆu��i%��#[1��cÓ�U$]z���������?3�9�)3c��3�۴�VS�&JY4��Y��-���5�W	4�����|L8 �&��}^`AN$CuA+r�}���p0n�{C�V3���gȰGc&I N�܏n`a�X:�,x0���Bdv�Is]>�m��-�s����;7o���v�K�GLoo��>�l:��3:�_ф,��V[Fɘ�%����c;��� 9�s��矧�3�����)��Ll� ?��/��%a̯�@H�Q,��u�ݑ�ޤ�Ƙ��&�D��
���+�:X�����~AF�8�D3�mkm�1 T؏��sӫ�� ����K�?���s00�r��)�.`@Rjp����'Йg�q�e��++���j�_Aޘ^�O&o�c�9�3��|��5o�B=.��R.�h"&6��sM��:cτ,� ٙ�*m��)D5ǆ�a��X����A���� BOD��$pT�R`�3�^���XD� N��,��rܗ�ZU_ #L���hL�[�� ���0�H^&vBdiM_c�y�e�� ���Ŵwt��2������^�ā4o�O.ǆÏi���U���駟��M�6���?�1k���>BV!̀j*Q/*g�`���I���:�p�13�@�q�2Ϭ��\p��Ll>�#8��6��:r_�:�~i�@3`?�9��i�g��+Z閛�<������`b���J���H0Yi�D��Ll.��.���\�t���Ϛ�B�1Vk)� �� 2��v������4������1Y�K�`�\oy������K>B����i��	*��+��2�lL��(�������s=��#��3�𠁾.�BK���Иݏ-D�k����(	��	w������
QS�Aޅ�c����'xtvvRWW?3�T+��m��l2�/ V��q^�<c�`���n*��577���A���
�
T��:�jŞ�,�6��B�D5��� �]�Sle��b���� �׿��t��1� ��7 3�Cc�lL��f�z3��_�F��O|��W����vU��b%��g����>�d�V��h=!�����x��)��S1)���	c$���>F�s��nP�s 0�}��4ɏ����+M��"�� `�Ű��}1Y����6���e�r�,����`�f�H��xt0�ƻK>B��$�aM΅U��,�м��U�"oz푓)�<��s���A���3t��6��J�``c}f�?�{�[O���dŊ< h�7&��npq]�D�/��X�/3�6�����.��c�\:q2=J��^&��Ll�^6n�� ��u`��^C���l��V�sAF�Z��f�gp��04Box��f)�Ѥf�q����㨶�Kry5χl�xGbѵ ��_����Yg�E���O�^�0}�h�qd�$�,���J�?rK ���?�)���	M�v�e�H̲1�?�3q�Y�2�$NU�����Ve�RD�B:�
���K���62�'W�xC%cu����Ǫ9�"Kۦ�����0�{������D���	����p���ԋ�`{VʐBM,ְ��wv4ۢtf2~3
T�P���_EB,�)�Q��L
2����S ��q3r1�Uo�����6����Jo9i��%�@�"�5y�Ɂ�j���׬�y*܆6&A���K8��?��pn�3�Hʾ� Hh�-�⬛Q���{BR-�kf`R	�}uu�Z�R�( �̽un��1R`�i�d����Yc��$�a6G�GK�2�L��PB����XJ��Yu�T�y2�L�[qΟ-��XB�ä��"Bb�H��<}���[H�k�,�����N>�d:���=���?��F�@�qv� ��p�����[��V�l�2Z�f���)1��^��"�2�Foe��I`N�}����u���2�
����i����	U�]�}�I ���a�����0�X3�Ϡ���"�9.����@r;
"^�m`��H�2��\V�"�D��^�**C��ғ���۱ m���R�[�⚦¥�n�\�R��X�0k֬�n�o>�x��wM�v}�hQG�cL�`�`3���dy�'�x��bŊ��_�2ǩ��on��"�2���o��O�)�����d81ȸ@��C��&~��E����X��@̘�qoãP`��H�UU 8a_�d����b(6�`�� �	��,,̲���� PE�ߌ#&� ��7����j���Z�Ӌ�,�/�!��t�ϸ������� �8��TG�3��6�n/ލ���z��;O���O�m���� `�yL�2���R)��4�����}�k<� 2*�yU�N3�f	Wcf+���^"/m�j_�Aŕ�~֡S%�}��nX�������+� tr�[����WqH�����L���d�`.%\��jO��d�Wܡ�1����K�F%c���XN���Z�4�]�U�, ���2�tc|U+�4�= 9f���ѯӲ �E�V�5��L�a�J�%�b ���M�c3���ibYن������ɿ��;�L7�t�p�皾M�4����U.�V٘��2�U?��]��'�q�?��ڦt�"�%�W���XODP����[Bh��17@ �ϥ}jb�e�B�*p�#�5.[ EaXM$���V�# �aAx1�{U���7oNCŖ�f"�i>n�*ˡԼ`�3S�O���2��S���`d���6�� D��Є4�j��Ȫ�� ��ϧ�,3���}���95�����.֮]Gs��K�5��0o-kڃ��?���W�r��+��[���W�{�y`�����dVjwf�Ɨ���>:�q�MD�2�f���DB�-b�%�YH�Oj\��
��fŤ��fr�l�2/ȅ�T�$-(�b�a6k��i�1��3���&
���]bp�0o`��8��<��q�N��
"R�YL7���y��-�.�Y��ɳ�,w����N�2����4c�t:�3���Ӓ���.D6l܂
6��w_�G?�Q�sޛ2���/�"YZ^��u�cY����ԓ,��&Sm�f�I��6���:<l��<�W�1��Ntb��df!�"F1qSS��3^��'����aL01F��P�U� � o��a���������<�
ѠN<% G� �����	�:�X�!���H}�U�|�q��G?�Q��Ζ���������4��=��}����W_}�+_az3lʴ�f��4�TNށh!�SQb��i�� �i�ػA����RI��^���9�X�%#��o�/&Կ�b1��4�An[��M��@7	��fA�=��W�$��l(��xN��`>O|�{�� �Tmo�� 4 ��m;n�%Aã^�V`��LU�U��"�To�����|��x<�V���DWc,�bK��Ph�+ӄ������>�V��,[�^W�`��4��Ւ)�Px�1��\@M765F�V��%���LD��'W(�)o)A�Z�ݰ����b�6^@�/�q����^xa����+s;�N�zΐu����� ����: �m�@�P�P��Bx\� 2I����bY����FIGw/� 5L��k���!�@��U�*���H�6��%�X�<�rTDSkn�u�I��l*:
�s��Ҿ=҅�����H�մ[Z��ᜡ�	�~�z�o���?����{�M�ҵ�m�Tf��.����W6�AF-�����g�}�Fx4 �h�tf Jډ�Z��7��C|U�e�0�8����y�㖷6V�}m<K�� ����XB/q���KV(E�"��z�,_��;�A[3ë,?��L�M恕4�FI%�eb�D*��K�~E��{0�����0U����@YAC���`z.��{�(d�$��� ��R� ��/~�0g���t����2�6Q@��	�֮]�ǟ�qW,sB1k/�`�$X�Ɋ-o�u&0�D*x'P��Ɵ1���"�
Ty�EoB�K
IK)�Q�Ri�z�D�N~N�W�h��{܏��$򸕅������]0��R�XJ���^*��u{�r.��ըWS�Q`��LMd-M��`"ӂ��a��=��̆�Z兒Aj� sӗ�D���s-�`0��/%��i)Md�( �wZ���g�}���N�3gk7�V�X�7D���|$䐘����2�'� �hn�l����<�pG mV$��B�� ����Ja�q���9w5�+'rO�}��k�1I9�@:�F�m�[�}^'YO'��G�<KY�f�e�kiBxY C)J,�4\O4Қ�l F��	�c0l掯D�.6f���1檀�$�SB�@��ȚQ��ŮRG�����L�:5������C6�6����,�E�ؘʽ�edR{��_�\��[7?���)�IM�������
4ی'�j��|��Q���y"1�U�y��LjHțI.�$\���;�ޣq6ˠ��v؛u��R�A`���R����In�W]8!�P� �j���-"�ܸKDiǪ�
����h�9N�+����7�,j)�V"& -m�2��Y��<��h���O���a����bjN�$�'�M8��-^�8��w�]r�%����s|T���D�0�͑ͽx\�o=�&�Dqsr��޿G��Ya��b�-7J�6�����!ao���J~�a�%`�-C^Ǿ���Л��0���#�����,�0m�\�Y��t�4I�L(�������r�G
e���R �K�Q&^b<@o[����ō/9NR�_�K ��O?C/��Et�Eщ�r���kw��4��V�x@�j{��ߗ,)�c��c�=���W��\v�e��r��V>%�W� ��&gB�KKXW�Fa�V�q��)̙4Ma�Ƙ�%v|���o�?OA�ř&�Z�d8�Z�'�;��WD2!�ތ�2i-AM;iX� M�M�:L3��S�}1�A���
0��t�~�U&VSx�H�k�Ńg���mcZ�~=o�|�
z�)o��Q��s6f;yu�}��6�P6QA���#���YQ{���ڵki��nݺ��0��K��yuX�:��Ic�I�RI��hx/%U
H�<��mU�,��V�ރ��b�3�,��K�5	.D�
�`@�g)��z3�\�.`����4[�b�]L����n���M���\���R�d�k}&l�>5Un�a;iF�Ms��E*�5,ƊBGaeZs ��� 8Y2N�چ�)�z~�@�ے��G�����M�6���߯�w�v�;�%Ιy4����8}��]��֕��yB�̼y�[�j��O>�䱷�r�^��%����b�{�ǂA����/H��2�ޘ�[B\�j��K���U:h���t�W�ضX���]��~��~��#H(�<��ǿ���Z^$O���0)K�E���R�Y��H_���A��������m8S�Q0P�J[a^lI �$�0u<s�i�
�*k١��L$���2���ی�W��z��]��s����誫���N����C�x��49j&4�� 4x���>�|�3���s�o���;ˠ��3\��{i�[ ��q/"n��}�*��NE�����I `�ю���*��#�8���+)�!��Ss3}�ʹ9�xԜQ�B�
�p0���o <�[^�3��uЂ��I��p�-qz0i�M,3���6[b��a۩W�T�	`X�P�.�Y�R|�8t�T��}$�}[OD0V� (#���GZZ���s#L[K}��g�كJɝ��|zE���[,?�p���眕e��3��^ڄ�K/����.�|�ӟ�n��hh�({��S_�p(A�z��*	���>^�+��r�A�楪�qw՘*��FƋԧ 䅉����'N~��(�
���G�13B�W��M��|��/K�L�1]�UVQ@�!��A_�k�Ώ���(�,r 
�`)9O�RĪ�bq�c6u��*�C���۫d6Ӯ;��,�SO?� �̓g�/�i�ռ��; �1�56�6i@�X���/o:��+����X�a��37GgM�5�l|/�u��:�Z?�Y��rZdxf�VQ��]��~2+S�dc������K�ނ~4��oK[��ܕ�x�e+���Æ�m1�Jѳ)�1� ��4���ԃVq;W�PR��啪�o@�]�f����x+�4ÿ��e�)�唅H`�m��q�R�����X0�-����I$������!(��E�0=.F�����,�ޝ�Nj �dS1'�<�ܚ�4����/�M�:��VZ��d�N_��hy�_u�(�{�6sO�7/��m�dp!1F�|��_m:��s+7�|3ǕAo�����o&�tP��-�X�J�g�.�+��s>I�g4���L1wY�`��Vd�����&��x$Ab��Xb��N�̈�5 �YbV�ȼ�b����B6+7�9\�M����f��p� RqO��B�:sr ���>;̑���wEa�8�|��^P����J��ǟHi*��|�`E.�R�m�r1x��:��6�骫���oyk��E�\0S�����$�� 2�� ��kS�c�u�]��]�J�s��3w{jno�6��$�b�L�mo9�i��RBh�FG������	\�}��Y�j좮���Y@��L���I>>NB��K�n�89�|}�Ea��y3j<A�ʭV���1��� O"�f.�4� U��~��L���4 58jg$�9��C	�ق�H ����_��X$�	O���9qH	5�X�pؓ+��� #�c�omk�B��v�y>�tӗ�5G�r}n3[B�&%�4�� 20�੪ߍ7��~��	ڞ�O�BӦMK]~�Il��]�h����P��h��ة�����nP�9���Q)��&�寽'�2�]�&υe܏x7�\����d�əV���+_���a�s�W�
��m�fw�,�� D|	���Y,ze��ɴ�&smp�YB[�
`��>B�T�Y$����(�p�5��(�\ 8���cz$�*�BK �+ؗ���
����Z_{��c�����rY@��X�p����#���_�b��_��Y��j���Mެ�VP��?��{���
ⲑ� �&}�Zjs7�\��ط� ����'��g��h��Oe�S��{�}N�I�Y�wN�Ҙ5|Þ&<�6��hV�XQ��ar�o�ٔ��a\ݎ�5��-��"�2K��x;U?zT�)k�L� �nF�3���$	���D�$�M�3�{�&�������M��_�����aUt���
1s,�N3�^�.����Nd}������X���twuӦ������O|�t�y��_x!Uo=ۆ�x��+o�*߸��QpA�	X�k,����0C��2�l[\Z��k������w�%�p�쩧�b�)7��@�y�\ôP�/c�3�H9M��۰*�ę�a2_�g�p����pX������ ����<�\y)��#@�{ֶ�8���Q��U�zU�R�
g6�4�7���t:�+��i�^X�/�L9�b�i�1 �� 5L�dL�,��r��s������KCfM�������:;i��u<��x�1t�W�޾Ǵ��.r.�^{�Ct?
�M&�a3 �;_��̣��O�Y�е�^}�������w�ջZ�&�hH� �b�9���M6�J��G��߶:��l-z�WW�LN�p�6C��վ�u t+�Y�|	@'P<�4޸���gi�$�l� C��iFC�G��Vz����r��f�]%�����2��ǣ�O�k0���;Q(]	-E9��˿E���[�i(5��쾦tl`4T��߁U�������?���͞;s�WP��%��v5:l*�m����7����9�Yy�J�_�F�l�2z~�Z�84�c�@�Zf��m�ġ�"� J2�ȣ�P��tg���>U$�.1c�
�E��ט��hHճB�^�w]xN�3�̈́��p��iٍ�?x���`@��* ���"��j=��Р@$���fF�ně���L��cK+�%��ŕ��>k�1)VM��Bh�h���t�;���c�赥���SO>M��2��]�k�����]7�]x!�?��z���n�bp�c�d�n�r4���z�w�]w%�#t�?��3g�`���J@��ָd�I��Ƕ��w�IMvQx�"O~!Ҡ
_���`!��hP@3y,�چq��P�X�X`kF��d�I,�"[��l+�S�Gb����� T{z���m{ԛ}��m¥�  (���T�7������o�ԺE7�k=�Q#Hl7'�L����d<����J$Ė�D�ڄ����a �&�n�6Tf���� J-B]�f��v�G_|1}�k�	6u-]���o�a��D��M6��%�sa=y�&��7<�@�/�>�|������ʗi�-�Z�1&I�R'c?]����h�Я�uF��i��VG{��ʵS�-˃�'*����|fƩR�z0Vs/`p`���v�gB�H��N�=�9$��go*L���o�a0eZ�bQ��^.I�����*;�y�J\۪Y�T�@ʕ�nO��z3�В08.� 5�G�u<4VF���$>T^&��[������t��I�r(op�=�.*l�6A�5�lj�{���6����8s�W��U�>}utL��ba�y�+��iDY����6���p!��\w^�a�@{������B�	<�J�
⊚Za�P'k6�m�ތe<&�j�6�c�Qū0�>-Ь�
w���p�ݮ�"�B]�sI�:��}�6͎�j2�h{�8e�l\1Ȅ���Ӫ�V-��ks�9��կ�,F�lj(<^��r=�j�_�����E�^{-�Ǟ�×���ﾛ��b�7$�� �9�m��L3���L��n��/h{�y�v}������X����b��v0��Kh�����U%���aQqM%�Ҥ��T
��.�g�C9g/E���1e7�3e�q�zތ�
�7q8�K�˛μX%�PwO��d�g�I��AKi��m�6���tf2��o�����Fi��l�L�Os;��Dq�$Q��I8���6V��Kcb�X�c�I+�K�� �!@�1{\�J��ΛCozӛ�c�ص�?�"����Sg0C��2y��ʽ+{����*�n�ч[Z�/|��0"O��AooH�֭��ӧ�@
�pq�#�C�;o�����3�.K��_C�
�L �r�Db3��Jv0�'%���&�)�4*ƍ��I��Ĭ��kF��Z�ȼ���4 ,��D1<�A<�=;p[�o�:3���  *��˴�&����+�<�/� ��e2orI 3��$�SO&�J}�^X&��
������})f�\I��O5�7�/���M�Ȁ����	!n|��v���t���o�_��ν��l5��7T�0l2�L�j����z5Y����ܖ�_}Mϧ>�)��?�6�u��@����Ji��P�t)��v҄��gUb[Xʴ�G��H)��RT�+۴���jƫ��k���x�� ,IB��~�E���jXVJg��g�N�r,%�
xr��̔z�,=YZxu�Sf����c�"I�5c�d^�a��� ��a*v��^bgP�h��'bM@s.�����~s�U�^��y�~�94eJ;m�Lh��멹%���j��C~�p��
�Mv�\`��Fo�
~�`A��O~��⌞4hT�����`���ƪU�'�#1Ȓ,q�vJ�9Y}���xf�@�]DKɱT�[M���(D7ǿ�
@�;���Ry���� +m��gzق�r�����3̊	=V}���6���d�t�TrA�g�H��!��o���X��m���oƝs��8V?�U��eA�T���	875�<�� n��s#����3Π�>r�w��n�q\I��Π��S�� ���d�����3w�u�A��|��U,Z��������?�-����$���$2D1X�����u�VS�V31T#3��j/඼��Xn��S�u��>t��/�e�/5/��7�j��r�<�@�}CgI`�8���U0� <�0L��ȵ���Ɛ���fmmm���8�v�H�(����dA�iY�hh�{���^{�pq%v�@���9��λҥ��N9���)�|��	��t��իW�~���N���na���
2��emִJ�]˳�N��k�c��oJ���j4��wؑ�M��	J��q5d�1VuP�
Ņ@���X�ޮ9�W�R�����&����j���zxYj)�>$�>�$���ȴ��~+l�X]H�S�%K�$l)H�|�p��3��׊o�E�s&����+�*J��:s�L�ꍬ��#�1
(�o� 	��b+�/��6 Ľ�ڙ��f�a?.�2V���55�v���zn��%,��Ϛ���b���JZ��	�l2���+8�.[vy�xl�
��������������6�+" ò�
2ó%˚����n������������q[��;̷�2�PQ^%�v��\Jz����f7v@ڕ,��	���k�T*K�N#�&�0'g߅�?�B�����J3�{QYnY�q�W��[=���lH1�Mb�+wwu� �ɼE�dT� HoJ0�jԟ��3��<c�ãqgp/..����
q�k�������h�A!��w�O'�x"]��Kh��� �	ͭh�l��uU�띿!�����|���{{�1x�͜e� `��G��$� �^Ni�>������k�k��/��������xL4�'�%�E�&�jg��»��m#�$}��?k����&#F?/zB�K�L��Ѿ3�Af��@4�p��{[�s$j �@�2�bx�BC�f��x����--��m�[��(�!�E`GG-Z���e�O~bi��vmx�m:�e}	
� �%v��=��_4�~{���^H+�{�zιg[*�ƍ�:�M��"�P'�:F�t6L����:Vf��gom*��F�u�%r9�	^Fu=��Ə�@�۬hd�8@�t^�D"+3*��<��(NC`�Q%�֖�k&- :JO֐ӔÐ���i�������WN�l_���f�紃�ij;Y���@7���V��N��/���#N\�����,��
y2��b� ���O=u��z�V���R��_�"��?H�����5ϙU�ޜo�{����G`�nm�K6�5�.s"��Va�5��A�˱(n�(�lgE ��o�M��$�f%8`3�X����F��[������n?��Z2���͉2R��ت%G*��vr$�8d��f��`UĬɊ=l�  Y�%ò3V��% 	Z�����f�̙\g����:Y�i�MwY�G�al؍�GӧL�P[5���/�}jk��DՓ�}�Zf|�skVS����|?��×ЛO<���?h}|��E/6��R�5K��W{f�{r�T�p\�v�V�̖Y:-,���JZ�9��?��������?C7�p=��'i���]3��_*�CJ��Ұ&����~��
����~�RTB�÷�t
6��i e��X�W�Pa;��ȀMa�oi/f��8C�V��'�}+=�WU��I^�
 <qZd4�KF��Y� �^�7�s�0|�f�S��0@�{s���܃l�o|���ދ��LD(��� :�>��6wn�Y3f�{��:���E�-08����Xn�6S"b�Tؠ� �a� ��ޞ���|ŧ�=������'����6j7�;�kr����+,ہ�g���Qg9���`j���p
�T_�ͅ��7��U<IZ�Y��x4P�.A\boa�(l�v�d���-�'7��V����
K��`����d�J��EIU�+���b ar�Ugּ����Z��[����\"�Ǽ�{��s�%��"�
�ń�o�633�|�+��Υ��í���t3�=y'��|+-�ҭ�%Ƌ)n�Q�d�o�F�n�WsՇV�o��:�w�������mJ{:�97�[���Cvœz@�zT���È���p?xۅSUh}3i�皐��I:����*�6v��ME��P$j x#�$T�D�ȲΒX��P�%�u����C޶*�0[��H{)�d�2��j�JR�/�����`EI�Z[�z�{l.�ӦlB�,5�v%㨫k35�[h޼�4c�Lz�k�K.����s�c������4�̀K���z�`F�
��2k4�z�u���^�������SOM���/�/�{j�P�N{v��<��f!A�K*1����`0{f2��5�m�JV��k $�*a:�X"��D5�ގ?L��85�T�cR�.%��֞4�+Yo�0��D4�E
7���-'"����z�����v?�H�[�J�`������D��VQ�h7KP��¥��ď͛7Swg'9�t�,c,�``kab�^�q'փ��p!]r�%����Ҽ�O��?_�W���k�i���.7�b�G�-����s̚�}I+@f�ϩ� ��裏&��?����z�jZ�` q@���[���z{D 3���hdi�����'M�jx�X�&�ښV�����^��B�J����
S�x3�\?����<�I�K+�ݥ.+Ȯ1&z�� ���l�[? �3@����1Ͼ���������iGes��ĪL�Y�����J7���ҢE���sϣ;���֓N>�r��g��6Z�_b<�1��XV���X�n������|��o6^͆^�h��j�k�o �Р �`H��O����ک�N>���z���!j;��iH"�*��XSSQ�4��2'�6}}�d�Y��̛I"KGF� M�'9o&ͽ�������h�s�LM�~ �]�7Y�����z��w�V�K���|�JO�=���V��JËҢKn��@:=_�hJ�4:��o�.��v�c�g��^���ߠ4Wڗ	;zY�*+@ft>�OY��ҋ.��n��=�^��W��x>�u.�� ��l��ܳ��*5K2��3� �ql��U);N��ڛ¶�yB���9�&�B�� ��A�9��4���5E���tws!&�fT	�)���6�͛S�fqi�U[]0=��lG��C+;��K����}���-�n?����y�5�:�+��uQ�?F� �ѱ�������/��unSS��͛l�2��޳�����V��y$�4_+޴�mw����+_�{�$*/@*Y��fT1�,)ԀM�Q��GsiêTȳ�w��tZ���\9 ��k��>?LO���7\K��
I�|��@��G�L�}/V��\S#���2�Je�(A����/a�HZ,�S���W[
���i~�w�{�� ѦM����SH��s>��9��d<��6q�͵�]MGuT���W}ù������>-��l�
��.[f�q�o~ߣ��,�¶� 3:���Xi1	�G;������Œ�I��$��*��V�ftTR���v�(�*��f�Ii��/�$�6��BK$`�����G����r���b:1g���'N�/g[&��q]h�?�@�����V,�5����Y��2�+�'��20��hm�2�XXS�����̸�]"��As�iS:��K?� C2�����Î���b���{l,Y2�c)Z�}��s�9����o��ٴf�jj��r1���ܘ��{nȇȶ㔜M�8��'�x6�R�-��(s�+Y���*5T��wg=njz|�����$4��7}��&fN��"���^��	�j~OC����x����\��P�#��XU�X��U^�����\����}����,�lYG�X^��,����I &��J70L���ƙ؁�g�J��&Ð`0L.�g�C�N	�A�B�1A`cd��"��-��rt�������N�Y��������{�^ԧ��߻s�5�|}����jA���&�2���А����q�3�C�u�H�+��o�w���*��C��+^A�g��얗\������;#m�}`W&����;QT� 2�������<��7�EjM��{&���u�� �$vòQ�<��˒݊��� �P�p����J��q���W����z�P^�	Y�D�'���,���D���6,Km�)c����D�����(�{o��!�Z
��^�G�LhZ�;7��$]�~Щ 3�_)S0��#C��o�{Q���I��L3[7��/OOM��pl��i�5Å�,.�����#@��&�okL��������O���]��Tc���
5;���w�]fܪ�K<;a�1������7��������$��j�du�����倯w�.���;Jj������
g[�f\W�ِ G�R��oV����iԠ�OL\{�ܜu?v�e�d&�֮��U�XR�RX��
<�>/9r�hA��h�"O����UA,Nh\*�{�0�x�;�Ő�6����`�}�����I�b�NZ��v���R���%ɟ�p�鸻D�s��u���8G���\����zM7N `W[,��Ņ�d��fȚ�7\�M)��s�$���f᪸��(�^�X��"��[���3�����Q��1�۽�=����@dzG��>�Y:���Fd,�u-y�g��/�E"ْ����i��<1���f��2Ӳϻ����\2.���X>ɕ�g+ѹP0�T㓻��h���}��皴��i�u�<��oG��/Q�T�a�D�sn����}7�ֈ9I�Aa�B�ٿG4̣��5���B&Җ��%�r�o����&1�3yJ �o444,�'	�H�FSą�[�LK+�<sI��{���q�v_�ҕa�`@dz ��yۧ�6���y�m�u����l2�KV��Xx�>��1t>���1��_�%|VK���yji����C�o�9&�u�%�6�Ɇ��'�]�S�;Kdl6��x��t����M�v�l�$����\ׅ;9=rV�h}"����ZP,0�\�N�C�^�x���k�-�����"�}�DX��8Arn3�њi�xg�z�����]I��������|�I���?��v~�r�J D�G|�?Kw�qU�Yd	��F�*�S-��L�ʪs�tvC/��D�q�-�}���n��R�-��jD�̵QRٝ��]f�U�g�*.�-�\�'n���F�*��4�AXo����d���}�8��f�w6+@AB���ݿ!��ʹ���EŌ��vuPY*�1e��ˈ�lֿ3�ed������YMųIcIZ3l�pF��6KGp�4�\�N�9iA��kݸ��P��{�h秤;�����#L�����������dg�\=vM���z�<՚�!��բ9)�}�p��f;ت0^�ˁ-�����:����t8���J&��6�ⱹ���-w��O�cZ"0n����d���VR~}���N���v�Z�y��f�Yһ���{��̓I����P-�ٮ:��ת1�l��)f4�wA�`��g���mf�v���ˌK*v[z�¥X�3.�49��}��u455mb9���Nɢ�d�f�W�$tAK.����0���_��mð%�ƮRv��L���uZL\�ov�q���ju�j��h�Md ��OS����)&���_������>5�m���K��fr�&g����*���2*���*�<`���*>S��z�M7I�2im>=��%�XM,[o�<��	�˻~�P�������� 1A9I&�|�'�Y+�Lz��j#�	Xt�hN|6q"E��Լ"ǉ�1_݉d~�K����Wq��}�B�P`]^��D�Lf= gP�+�l��ߥ"�f�3	Uʾ"�ex�,+n���9/Ө�c;U_[�A��6�;f'�	g�q�L��_�*�4��Oؔy1�����D�_��� }���_�.�(&�<�3]�O�޽��;��~��&�4j;i�\o���E�'���	}i_-]��k`�d��ºB�V��u�����Ko=�%�Ȓ?/��F���G�<�Id�3���f�f��+iW�u�Y�I>mo��ʈ�{mV��,�b�oU]�D��'I".����EM�l�&���t@Q���+��1�@U�ݑ�F����`�GUp��}r֜��r��N��NhXX�9��k��/ۺ������z�G��O����Tv�FK�����L\ye���&��U���DO=uT[�M���iY�[k��MEU�R�F���Z�dw��|��D�q��f����J�^�����ሞMb�;������LZ�$b��o�l�c���w���8}:���}G�,�(�$�Ykm�_l���B�9^�|���ɟ����N��<m9T�ɒ���%D�em��<n
/�"�ӕ��r�5;>�8�viv"°�x՚X7Κ��G�E������Ƿ�w?p���69`\��Yz��|t�r"�7����k.ݲy�7��M�`kRu�N'ON� �*��r�[e�Ҿ#s�a_wˮ��(�T��e�M�3}��6X������-4.4�9�����G6�/��{P�,��-Ԏ�K�R��:Wsc��t��db,I7^0k;v���+��G��8�����	=l#J�2��%CP��$�S��Veh��vu�`�7�����'�M�9�X[K*��B���Է3!h�\2�Jb3H��V�D�?00(���s�2��e,�>�5c��"���i�=K^ǯ�4r�k}�|�!��?�S�k���C'h.��b�+�D&�μ-�w���������Z7�5Xl����y	ڞ�l`}�����S�+I��)8�l�Ftu��"�ྡ��5Ў���Y*L4���$�2�^�p3�7���duY��ڹѲ.�0����,�����JV�^pn�F4/Ѣ����z�1�Oh9e}V��%�@�t��X=uHfZ��%��A%��^��^��t�$l�%�	.k׮�����rjzJ,�֌ͬ��O���w<��3�������D{��j	r"��vU骯��n�Xw;N
�`rx۾�ei%�����b���;�_�Z���0Β�۞��w�ohOCO�#�}�r�riN$C������Q[e�yRH颿x���r��>�S���I��O/]Dx��)$/e���=g�=?�=a���;�7�Ť�T�%h�:1V;��b^�y�������E�Z�X(�jԖ?[$I�a�q�"4#kE\�C��b������
6O?�$�ٟ��΢��h8N�-�e�No��������k���~�̌����y	l�C�kF(~nq{���\C�76>x�rߝH&N�l�:wr;�3R�ov
o<�ʋ�I�q%3=1��J�b����~�YŊ|�NE���BȦ%w"�b�gKʱM'�Qֺ�=�&���9IƔ<�Y$�-�#����R���^h	�q�|�I��KId��'�T뵴+R�M~�)�T&��Z����0��g�4����U3.;)(��^}��B�����߻����Ƀ�{����5�o|S�?Ed5!��~��9���@9��5�Kr���&�I���>U�Z\&���~����7�Ѹ$�����~;}��K�ر�i��Y�[�O 33S��=�vȌb��U�����olJ���bc!J�؏�-�Չ$��I7Y:���z2.ú;��b*�2�%g[|�\¾oTɈ�,�q�gI�/�]�x��{��]��8�"���u��q�L�o��-��J'D��l,�(��yq�KQ���Q�~�J��r�s��y�w�扔֠��ߙ��*'�����,���J����&,Ӷ�����t��qٟ�q�jXd��Ӌ-Zl��?Ms,��~�Ԗ��ݻ��[���ϼ\��^$��ŝ��;��d��H�&�<x��!����RH�+;יYm��}�l��q�4��rQ�����?�>r�G�⋟k�+k��ޥO37�-����W������G�~D�Cr�s����O�g?����5)'~O�j����K�E��L����M(�8���St*���r޵D�hd�(�$���D�ƌ¬hd���ƟR����#��[�ɟ]Xdb"�6��v`�r=�m����曧�H4��K	�}΋?�	�|N(�Y�>W���f�!��Ru.Ҧ������������%�.l۲xp�f���p�4M;MSb3����<����[N3���7|��<~�o��K��W�>��
�D&��CN"�voصVtW�5��l�T+՚%9�0~�g3���2�[��J�����+/z���RCZ`xb�;�I��cr��/���;�S���9�#OȻm:�t����� �7.������X�"��u��⧚?��^�'vvӄ�=؋,	�� ��:���>�zm�����mI��$aQſk\������1�J%u�����I�_%�P*�Gݭmo6J���1B"�1�R��a�)n紟�&�f��Q��2n����s��4���T�����Xg�9�����__���߭V�A}�.���;g�I�J�|ϋ�M��T�7�liA�_��׽p���������3if�2k���Y�x�c�W���b�KmA�^e�"�@\� 29}0�L̜}"���\%y��Z���{4�W^�+��.:����oEeF_��p7"���_{�N����mt��?�_����Y�җ� ��Ǣ��T!]�w>Q��{-]�!~��J�{L1�<%��N�'G�vi���ŋ*�Th/%Hʮ���y�Ix��-)�����(u8�x6o�o�~�J��aR�͉�3�k�a���l\ڳ�H�<Zi�"��	1Z�FF� �4� T$�ٳ�ʒ�ㄆ{��v͌���6#c�hkf`J_&bkF�����B��^d�LLH7򑑵4q�8}�#��������� -�sz D&~��I�%H��9ڥ=ӄ1�y84Ezܷ)j�h��CV�^����
���̵퍦梋�K��ۿE/���)>kF��唽n�o:f΢'��ַH���'z�!��7�閛o�o��-��n�CURQ׎��7��/7���e��f�4�O�رc�d�Ēa1�¾v�Y���-�]�W�7�f��.�*�:��ǊP$F��b1�s��������[�z6�����x��0~Z�k>'��*��%�N^�	�U��s16���e"��ML����6j�����4U��ڊ�d���>[�{�Qi���M:8<(�.]`�`�,.M��l����UU�vx�̋iZ�X��{C�	�� q�k���ǳ�whnj�r�����&N��P�izd���I9n��6������c�W���Ɂۿ�z���tп��R�)��ڈ �zO��U���N�kQ��_�Bz�^��jo���6mV��֌���_���o=��SO]{�=��A~������=~�q9��	opͰ�4X��d�osLfÆ�ъޮ�+��Tvg���Q99E�ed�/>ɦ��=q�TAd֢���p��Ė��[��`�̇U���"��ڱ�˽_`!���(7�������O�I}����>��|�.��~�%/�/��~������O����������ȑ#�?��З�|3=v��L�d����V\��QDh�U��"���B��%c��ڥ��g��Q_[���U+4C�C4��?V(��m��(];a��}���������akE"�]Ŀ�YZǟ9�a�[O_ͺ��2Ř�V��KU\�Hw�9��n���I���}���ܙZ��>h��4}��Fߤo�Π����
��w����JE��z%�bs�}��?.V�8�5��j���&;M�p�R5jN}m�ެ[ڪf��O�駸�fvH�K�Ì{̝��.�L���X1��������+���	�	Y�Vܒ��d|2>y�I�x����7�
}����O/|�蜭[i������h˖Q�����:����QOк�����w����ə7Ӎ�ҽm޴�&��0H짒�}$&c[Ű5���i`p����ű�'h�C�%�����b�HfI�b����3�fPjg�������棆�J�K'�U�?�s�+�[��/A�f���� [1Ebݺ�����&��Xl�[�����N=u�p�O>9:��	��>��wQ���u&��͗�TR��?��A�;��~���?LO<�=���i!�&��~�<e�&�O���!Ia�l*n�@%EFى����q,�n%��([�.1����Mi�_)A�(2�_d*�9��TH�E����,��]v)�c�ɨ�З<���Izݺu"��f�"}�����"x�K_F�^z)��~n��M�b�V�7O$�6!�ԯ�u�+i[�sWޱ�}����;��:p�-Ri�1cD:���5#����*�e��g��ߢF�6��v���⚜�dkE��X3��9CSK��g�`��\�f�yƲ��ş����?��8{/�՝�陠@d���k�=і�K�@ÄO>�0����+��c�>xV�Z�D������)�\�?w'�N^6N��N(������9-]�'�GSJ�F�)��qI�z��������|W[9�����6���,<Sӧ���Ez|�q�^��'n��1�z��S�Ed�>�ha���=\3�P�Tj��ݕ���1ez>u2��~_��yQ+��[3���i�龳����<���A���V ��~��K�m���?�^����-�����!������=�EZQXX����*zI�*s��O�}h�G�u��_���Jڰ�?Ƣ��V@�Sm$Oii�߭՘��I�iV��H��*�%��N����ߝ�)6忩���ifMS?�����k��69��+������{�)�ḏ�⮻���x�m�.��c}�c�G���!���V��]w�u�~���K`�>a�Q��q�������gc5��'�|�\��=����?�������C�;p'��w~��:uJ~C�Ni�d
~�MU���]�Ai�]��y��=Y��!m-�;qw��Y8���u/f\�8�L>����	��ٔ��m%���q�މ��訸=/z�s%��͊��w��C�m����ᑐ�~{��ۃ�����ծ���7����������Ȁ�t/7���d���m�ݟ�e#��$,$3����kق���7������'���݌��]����O�}�ȟo�C���ӊn�A���J��t���8+����:%E�Bܐ:*�u@a�C��]}�Yg�E睿��HN��]]t�]L�����A7W�hg����K&��g�=�iA�g^3��CM�[�;p��o��G?�G}Dn��|��2���*�q���1�
����KLA%�I�ɖE��Z"n���Ӊ�k�c�f��m�ߕ"8I��s1m:s�ʦM��Jٺu+�x��Z���Q������$�}�:�_@�w/�#�z��Nڭ�D����m��K/�=j�VBck��J��TN����&�b����+���F�K�p8�l�
ǘ�o�1;I�N�}���bMv��v�&[.6�/�9�w��	.6�Vo��{�?���)� 2�!R�|P��*�#K=�-w��<�b!����k�mܭ�1F�6���.3�hX`Τ�p�vz}e�6-@M:�]M_�2�CS�y�s�x�����mݬg�/��U��O<EG�>JO=�M����S'D��~�i�����Y��;L&�&l9r<�{>QnٲE���,&|�q�F:��3�Y�z���d��A�N��z2�K�o翕I�3�c��#%DX�����m�w�<�e��hc�}�c��۷���	 �eg�`h�ƪ���6VR�5��&)/%�n�XkF��:�vG�����3��AپV3M4]:5�Q������?��?���������U��=�B� �D�;��r�Сȧ�U���&p��kX.�u9�_*����&3*.Q�/��4��wT������1���A3-�{�_#]V�r����Z�GU8p��
��"�"ĳI���>9��8����s�z��k7'��e��~�E��åm;����-:�!#M��K
H'�p;MO��{���{|������߾��;��E/�����`��J=�L�а��3��Ș�檈�w�v�B� iе����*ґ�3Sg�2��n�|�U�m�/ӯ�9�@���o?G���!z��d:a�wY� g1��%"�e8��]��v�5:)d�0Wk�\q�Z۶m�C_{�i�D�yD�}���}Yx���������u�xm7|��Z[1+�?��?<v�w�7a��	�
�n3����7L�^�g��;�O�l�^xz�Z#��4�h<c�h�Ђ%.5N�o��o�^x�c���mr����u��?q��[�۲�X�K 2]�c2sZ1�,����]�'�g���B1�)rIT:T�'���	.�@����p'�oYXX����P_'�H� !Q��I<���H��J��O9��K`��G[����/���"S[3@͖�,����\re���34S7����!��K3gr.��!Xd�}v���"㗵5â4�vXDkJV�1@�#C���u3ˆ�.�Ae`����������R�k��ݗ��^5@d��ؾ��7�U�:&k-�0�F�=�戩���p�m>[��RK?�8���O�n6�Lb��t������iG���V:�5�\�~�����ی�o&�έ_�R�ec,gq1}QkF�~ȧ(�f8��bJ�O.�\C�Ӄ�~l�Lj��4��q�|*�ߟ���U�����}��5�r���K�(q��Gcw�%]P���� 2��c/R�ﲛ2^�e�k��f�\Q�J:I�W�ɗ�ߧ�.�Lh�p����~�\1��C��J�v��Ǣ�U˧��Zw�$�y"�oy˛i��ɷuJ|���lY�p"3Ә�"�����v�Xp�4��+n=�ZI#P��os֝�T
L*�m$�3Ф�L�3��e҆�Jw��C���<�٣��+kZ`�y��;cګ"��;��W���JV����~��*r��7V0C���w�uǎ�O�S�4n�h��ә���פV�%�ѧ_���Z�3-��̯�K1����f0�e�o��2~o��YfQ�@��x�~����ylt��f���L_�m�;��Zl_�vH�)2ݜ]k�X-��Rm�ͺF�E����d>+"�_��e��n�߹�zr"�A��LCͪ���Ռ��]��4-.<��orcX��fԥ��[Nw�k�e�~�!7of���ς�?{Ɗ��Ȉ\�LN�x�O���v�>�-�*3�:�ި��, 2!��r9�0�d��:O<�5m&;r ���������ڥ/�����wʌ���B9��X\lo��t]Z��Xdl�n��T���
Um+׾H�n���f8&3e�5ܜ�ff����pO<%��������<xb4>�q0�" 29�=�'�P���.��p��U"�����8�34��")��]U��b^�K�֦,(���1�9X������u��ō�:x�M����暨�ʎl��3ͬ/��Ӎ����k�x|��돔����޾1=C���PԻ�V�}���251)M3����Դ�q�YT�C������S�d.x3� ��b��Sƿ�f9@d�Lr��`���ЕR'fh���f�z�&�-Ùn|�=o� ��U��c��5ӧN7p[#�j�Ԍ�BK���i���֬IvY���t�6mwX4Z`�5,:��F2v��}c���cYHIƚg,� �R��b�կ~����F�@o����i�!�~���)�h7!�͛EW��L�T�H��W{�2��@�����+_w������=b�k\�ي�����gVL��c&I�6Z(������׉�*�&�[w_�3A4k��'�!�=z�����>~�ɿ=s�="�+���O��Z7��jc,[��eބ����k�3Π�+ŊAJ�Jc����wo�o�vM���#[W�X2�	�L��u<Ι��?���&df���q4(�Vc�a!I�DK}933�СCWP�ξR��R �Ƀl��S�ɰ�p@EU���,� �I܎��	�/�fٴO�7�q�@�tތ���]��p��FA� �pF�����Oe����I'�$?�|���7\���_{�=�2S65��l�7\��fE[S�����R�S3��9L v�y�ےƍAH��q4OMp�>s��\5cQyRw�|�YX�M,&��D��@d�@肝z5�&xϧ[ϞZ�(��=绳�K}^ر ��/���D�������F7_�������Ծ��?�6s�aF6W��bÖ[/��d\<R\f���c���c�b:ZH�[�(�tp�K_�2�_~p�.��At/�3��L/a7���|\����H5������PR\�*�UhтD��M?~��5�'cI�l����Ft�K�A�������[oM?'��rm�,y��ex��~̉��HJ3��і��-��S�44�ƌp��>eI<�b��<m�g��������#�8�� �S 2��S���ο���a�b�ɸ^�B�c)���=�[��_�%c\n�l�Q��˾�-��Cu�3�O|�>��y\&ߘtb��XkƍYhI�K3�,������1�V2I M
�8����7��� �-dl�׶&�ō��S�����Z="�Kx�,dR/9m_")Bsq�r6���]�m��j��s��7�0%3'-8A�%g�m���:���~���/��m۾/"�L&����T�S3�ܷ���ɖ��,�Z294�S���4>�����x�W�)�9 8{���0��q�������\��f��𯸪inwNq$F��~�\�� � ( ;Bڳ�߶g�W^}u��d��f��f,q!%_��րX)^�����w	0�����!� ㅞ��e�[=a�4 �I z��czD��T�i�'�em�q���V&4V	�O���/�p��v�e��cɸf�Pfp�!��) ���p�^�K�CqW�%S,[&�Ϯ�:'p\ƶ>
��8%253.�Y����pM����Ξ���"������$S�N��{/Ѯ]�C��^��@dr�ռp�q�p�l_�J�qb7�Ծ��F��eO��xA��kVy��Cתv$m`�� �p_��x� ��W[�9G� ~H�#�N���<`���%ÌkflW�������ea�-�Q3Fd*6Q��՘�sVL�^}J��c�>J��[ר�4�e�3 2="iʧ*�eV�P${���5�q[`}�2�eaӧ����J��+7e�6S�W�����1���v���T.�я�.��@�	?h�lG�K��FO��+ͪ\�Bd)��8��f�)��h�T�i���J�hܲ�8�Pf3�ū��$R�c�6�F^���nz��_=�l�R�r="�Cܪ��N6�X%����L��{L,��EU� B�"n���4��\	����8�W6l�@�{��L����ݮ)�7�l�Ll��Ƹ	z�q�֒qsix�w�IM��L�L��=7?�(������̱��ĉDg~��{D�x6�_fjp�ri�戨��/�~�ǌ�.�盾o�穓�Wn<5���2�L�ٹD�x�hio�������ᦔn�r�o�{�k�-eؚ��d�Y�&���,Ӿ$��0��՚�EJ�榔�q�q��\��ϰţ�fcJ^��Oбg�!�[ 2}¬�⌘ \�	��ڰ8q�������|�	� �9ښ	�ب��l��eZZS6 o����3�z�Y3a৺2��-�1JFf��\o�6n�nf!�!��~.[1''N�-��q���}��bk�b�<�K���/0�3���bg��1�W�-�5�f[/�y�xU&U�-,�5 �C��]$E�5�,${R��@r�׫/�M�2�fjހ9l�L7�.p�[.3�Ɣ�h��95~(����7��𮽌�C�߶�فeX��t�6�g�D��L7s�i��h���}Ev@"�%�A��XX�aHd��󸭛Q��o��?����6J\��ٶJ���ۺ��1�&3��	L�c!!��@d����z%Լ�t}MȪ*�eY
1%��bVa���[��F�N��1G-�,�w��O?�6���?�UUe΍�80}��T���BfR�c��.w	*Vd�{s`����s�7%N��B��~����p�O������ڵ�n�:-2�S+li���� 1��;��v8�ȸ�1��I����UB�pg�Vܝ�O��oY�?k��^��.v���K J�ؤ�Wd����A`F����Fn�\7ck��b�3zŨ�����|���G�yN]?� $ ɦͯ<�=��Oxw��$.;�ٹe;賸(���w�&G[��^���$�F�=���(3�ǋ����_��Ӓ^[��4����5�,�L����b�X�E/hm=�V����LFI����sGv3K߾���Ծ�df�D�[Atɼ"uo�,N;�	B�E 2��%��t��a>���L���/���ԅ��D�W��	D"fΌ/�.(�+yZ�KF�Gv�og�7���*�љ�k�-��Lw� ͖�-4�g���T��]��Iυ��d�RŌ��_I��@���]��6;)�D��� F��<'q�Q&six�l�'y�z����#��8G���Q2�u�}9)$�mi�.��]ѥ+�əv���xe�雾��E�T���H�4?�*zD�;�^ϱ�o�$ V;\+����K^\�̷�+���MF4��3�xh;2sv�+��_�j��uw �"�E8�_�
-�P���P�8�zzX��n?�LN?}c4߅��1.�Yf3�#��B�+�Qn8Y����H3[8^Rd�����o<��x|�2Ҝs�� Fx���t��NF�_�K_-��!Z��z��������d�?�j"��,9?�jY�Zi���H6��eY�;��Q�.�"�.���Wl�Ќ�]��֚�"%��Q%C���e��vN��r/��-�b>+���ql��[�Ӗ?�x���OoM�4o�xV�oki��&1�"�ܗ�A|t����\�Y� 3?a���m�;����&�.��g��˩�1cg�
�v�~XM��j�X&�f��9���/���S1gi	ǚ�0s�&]vcP������T��X��`�r��V�\�|��VEf�/I�?�f�q��i��gk�Sv�evB�:f������;�y���|�\E�c;�D����`�^\h+w]Kj���︒�R�e Y��<��1A����V�
CA�@d
D������P���X��؏-���y�)�PJ��c<(d�\1Jq,WId"�`<{Q�+��-*�,30��H�B�����*�2;�s��޶�Ǝ1��)	�ʵf�*D��YqI��:��@�['�6f�.�
me� Dfu�#�����tL�eJ{�tk�Tw o�i��L���@�L��v�-4	ڹҲ���z%'��u�e�G�3��@d� ЌWk�b�W/ˊ͙��:#�z�'e*dҬB��x
Lʍk�a��*�cҀrQP�Γ9�r.�t�b.��c+�?�eKՎB����xQ��;�.��\��{v�e �x8�j�Bgٸ6������ɱ⫪�$H6}��i|g�J�6���TЉ	�v��@p��@dV3
��2HwX�DS��uƲ��@d�,��ѩ� �'3*#Ld�!���@d
��I�q�nݦ�s���/XN�f/�$�Ŕ�]z�)<۞��Iߴ�5�63�$����Bj�Ē��v�мo�|��ح(�ۤ�.�"SR�вſN��c ���d
��2���L��varn��dx��⎍l��h鋪�DL�L����l�����k.K�H�N�` 8�O,�������LH���w+8W&��Y��/�vm8�g�V6��9�_n���
�y��㑘8k%�}����;�4�n��E隼]�A�X�e?�ZH,} "�g"�������Z)�)m�$7GO3P �.Y�4�sl@_�Ȭ"�Sqz)y���~����V�#M{Sz�����Wvs�J�5a�lJ��#��ل_���M"0�fB
 [�R�qkq������t3O���g\}"S8\����8��8K  F
5	��L��:/ρ�b���abXS��9�t�ӏؑ毶�  �D�`��`	��i6��[�/�u{�S %�*�D�\~����D��;�pxh��&�ǽ�B�Y��)WZ ���+�q����������n&�Ҝ�u��s��v�	�S��]d��A��H����2�x1#�y�������v�o�r��!�d;��z�G����~�=�?�#-5Ώ�mF��@d
�"b1abTD�]�.�BHZ �t����(��6��� 
��v2f��~n�y`�����m�y2�L`暛x���fc2nkV ����Ia�>�5��xy�Ma9x��;��h�	�@��4.���E3m�|�/ 2E$tn3w�����Yt�'�c��#M�t��̖h�z�k�$�4v�0�=2�}:Q�͓��<����.[��M~���Bly@dJ�b�@)Qs�C`�J�;/i��?��L�t�C��%����|l����q���y2� �>�Ba��2rί�y��g�1�'|o���`g��L?QNTs/Ă��g{��]�Z�B?1K=1/#�ٹӪX�zbv�h�y!D���T���-,T�׀�D�p���R�u^*�y�x�B�!.`e�),����d�S���h�A�Ie�f�$  � �*������"S�l�F�R�w�BQx7���`� ��M��&�\*���&���_�M 2�`�rsL���4��"�c �D� (�A�%��������]g��;1Kyv�N��+ɖ�Ǖ�ϛm�4v-�n�ᕡK�Ujm_r@ez<�n�D��yY:����-��a�F&�Z,�L��Gx�c��K��8f������t��x��RT7 Q���LG�qu/�u0�O�*��ȡ��]cx;�Y�&���|�<nkn�d�Y�jZ���_Y���t���x���� Ka1���Ф�Z��@d���KB�\w<��߿;r�&+���N������=�B�B2�G��!#3�=�"�<�Q����ܿ�y^��|��{}���~�u��|�0F;��E����9a���%��U��5E���Ƹ�%^�:�{y�6�L�}� ���҅�{�䠤Ñ�=������$y��0�'L����Dk�;�P?�a�hԻb���0�c<����OJcjQ�Ê��L�6!��Œ˲
W�Qp:X���R_�0si�.,*;����}緅N$fP��$��8d��aʶ�ާX3\�d=7XZw�����1��X�_N�6�c'�nc�%g�8���K��d9�7t,�/��D���W�,��x���R���� ʋ�>�=ku
_����[�f��_Yɨ���X=��_��5�>!�Ѫp.�p>{�I��u�n�kyf�r�Ș�uUul\��i_�l�@O-� ��\a��I�x�����
��	2{��Ѱ�r�� ��c�*�N�7�|,�ViQ0O�2�,�~1������
�-&VI6mZ�YFYP	�O��� �Mb��bn_4�4ǶI��x�����4�k�mkck�f\�}g97�r:��sfU�%-�SlL��ZW��L��s�w�יPVl~����̥+�˛Ah�j>��
�{�FVru�N��Ch[]}1��]�I 5������$��d�u��r{�8��cL�QW�
���h1~�K���2LMҦd��Q�g�ʹm��l*�W��z�Meq�:�|
�݂���BF̈́X�ɢ�d����S,���$�|�迥;+�'��M�tL?cP����=�\�<4��K8���q�{��=%�6�p�'�w�����:��{�`k��O��9)�����4!�R}�B����4h\=��N�R.�2�P�o�4:��G"�%��L�a�`��&E�1��3}V;��>�׳j����������A��ʕq�2�R�qgIuϧv�sY�
C���({3w�3�G����O�-x����Tx�xzn�>{��Yx?7�j�(��NPa��%�s_��dLkƀ��"|�羥M���M�d,m��<l����x���7~�<��P����jh��p���(s&4x���ͷ��>���J\%/��B�Ӡ����b��e�EY|�X�_g\��������-�S�!M�3�])�P%����ߚ��`�T�����vO����^g.--m���#�k:��X��*�|l?�Rw7_{pBcn��}�Q�5���[N�KZ���_��ּ�:ZX5ݨ��v��"�M�\��rb^��a��&�:���o��d�	p��O{G�"�=�2_Jſ��|ʞs��
Ϗ��g8EX�_<��Ul	��]����)�Q��E"H	$f�:oX����
�WRV���`w�g���w�*�]j�ʳ�2�\�l�k�.׿�@i�l�R���j��5<��JH`�����n��X@P4Z@C�]=@��P$�'�L����*K�2ۉ��[Gp/$�C&G|)?�������J�';�K_�wfњ��;2�DDn_����M���y�j�C2���N��� 7���b���K�v�T~Z���9��X^�K��Ф����ş1x�4Ԯv�I.���9K����:���8h������䡟?�����ݢ���d[X��3H8?ON�*,��l=nݳ:��Ҁ~�2j�Eu�7�����H{���1�MkmO��ѯ3&�15�k��%�/]���7��5'ءF�E΍u��k���-�~�}���x�����4�$ef�ڧB��~�xttùT���H��t�WT����nN.���Z�~��D�}�ư9sG�|����x���{�T	����E�>�������Ƭ��r�6Q����(�l0�\7�=�7���8�ȗp�b��|�+��{�$8"�ǥ��ͣ�����q�1���[e>���޺��۟�� jKH��]�L�u�}���9�M�u��kwo���5��F��[{��=�ą�ӷ�����)�O�Jn߼��X`�3�w�q��
X��f;%Hd?��r�"�.k�n�r����S�W�+W�Dd�̃�i��^�#j�>����܍-�^ARfӌS�I����{�n���x�>��).,%�K��M_����NE!�QYt[��/v�2�ڲ���
�'��|8_����W�sY#f�ړ��B!/\���^�qQ���V�̣\���HM���㪅~y+���ki>ՇCc:C?��׏w���WFtZHm'���l<���e܉岪��&���^�P�����R�)6u3�H"������'������WG�`0��-8���[�1.�ՄH����C�z����p��������J)�erI����v�ù�:"�#1�fϗ��{/��y�=OF�:��WQƎ�ZyS���QE��-�;)�*I�{)��dr*�-E�/���mm6-�3f��z�Hq;x�Adk&���@��!����
!;��P����q�X�V8a������]V}U��y�K(�t�|}�}�y��,�H�Z�$G}�G����E����Z���I���! E����x3�N�ϨdF���i��m�[B��Jl���S,���M�x'���?���r���$�������]��n��g}�߾A���KDDC �����������F�΅������"*L;5Jz����]u�2����M�f�f���I%u�5�
�Q]v>����{��z'��E�B����P�uj�r�J�xN���?����Q�c37Y��9Њ�]������]��ח�["���`�F�5oZn~�.���V�ܞ�#����Wγ�D���>zf"\Ϡm���;2�'���/�k�s���u������PU<�k��'��
����)
�sF,夯���?�H��~���p��|��K����ҫEa�{�fV������?�3�}�cXA$��Js����~e�r=5u@�ᄲY{E��oǎP���7��ji�u�i��ŀ���6�T�K�8ʿ���?zɠ�m�{���(ՏD���̄i�p����v#�U��5�wuh�
O�B����K*Yx�>2���]p�����WU��ԇ��^�K�r�	�
���`EuFমQ�O�Yh�S�*�4{�C�D�w�AK��������ԃZ�D�✃�6l_��#��R���0v���}��)���RO������bFt����BL�CA���P���s��%��*N�~֏����B�ªL��m���bGu�?��w��;�{�U#lv)<J,���x�Ki�>��k_
�vcn��I�C�V�(�����>�t�Y<(y�/�%�MOr�����!�+?�?��e�'���w6�VNN�Xh�n��;�#�Y�Q�WzS�ZM]�P�.c��2��c`VM]D�)O�>N�	���J���;���w�^Յ,v���n����s��p(zP�?3>��D,�r$�z�ov�Q����}�����긝�λm^{�p�"�� ��f�n0������T�Z���B�#5!��vsQ�.ꗮV0����;a#N��J5�?�h��D��Wz�M�5�B.s���t���kg�i�d��$d*��'�.ǧ@�:S[[M$L���.pJF����5�t�]���:�9I�W�˻�����.�-&r�X���x"QXsfu�ILf�>g������G��K�x���4�Q�/�E�A�n�"�!
F4j��G�� �]�����Tz����ݬ�7"��+��kxm�}�"�-+x	0c�/��M�g�:���I-��#��s|�~M�� �Lk��?��Y�h'�.���@?}1%	w"8p�xF9�)�1�k��p h P���`�=X��J��l�qi (�V�ƛŖ� �-���$��jry���l��e���B�s�����s��}�h3��9)3m�6���ay����;{���+1/��"��u�O�p�\H��3��^MK�(��Da@�(O-{۪� ��Hv~t���O�A��3��z5��i4�]33c`�)Q!�Jv���A�8
�`b @Nb. ����p�1rw��19��
��}r�̚!���͙��~Yl@��ݱU����l�c�	�0^R��̻�e:`��L�gu�+3�a~l6�&= �Bv� TtsD�UY�`������]�oQR:Ǻ�  �1�p�x&!�g��4 �1f�4�y ���u�����1 E`ptD���yE��9��o�	o��@0��v�N�������l�����4�1H!��`����?�����-����Q��F��7��n��b�=���������)�qj�?�E
v˙@@ii�p�)�,ޙ���"�ߌ�~�Ђ�T�"r�.���P�?(f/.� &�Y�=O� g"�׉�c��1����C���a�N������6�`����.�#Ɲ8F��`\� J��	i��d~8xCAv�:v��z}�e�u�3`�����z��>b�[_6fA�*V�Ž��!�a|[��>�0e��q�.������]���lz��%.s�)W�^lL|
��&��y^^Z��^&FHW�&h�;2���|�Ǫe�n��X�K%`�T���pƃ��X@F��`(� 7�b&�t�
e���/*�#L�l���ǈ��zLN}0`�>��T���GC#zO����u�a��/�����Ns�q_%Z�]��vRCM��t1��"�4��x�-P5����e�,aT�m�b��k�]C�cmW&*�{��������؂{�3Z0Cu@�k'}�)�iW1��H�"ǆ��9PU��b����LB�����p��?�qnc��`8˛�������͙���g���j��`�����`���Ɵ��3�"#�ϥ?�����.����F��Ko��+x��{c�����<cF��L�4���Hv2_TA5(��"��J�ށs�F�7�	�?�4ySC ���H��=2�<l�g`X�-�5�)ϱ�jc>O�G�ǯ�1A}䦟��`B#���QAz�<�e�Z=OK��k=	Dd@�Q��K�����3���rxy�5��tc"D�A��]X�b�	�6�_>�8=��_*��$��Am���]`xUTݼV�A�]��@�����s��_�qp�D�s9�h��i�����!ʃ�����& I`�s;���h�T�_NB�)��M�+{؀(T��Z�32���i5,.�߱���X��`����D��30�M�i�����ܟ�݆��uH+X��X�op�a���k
9U��WvM9eXwq�
>n�^�.	y���h��x������%�F@�JV�iә)p�B�ʷSb�vd�(;�>�d�b�ҷ4.��h-z��@?�}0c�@�XT��缹JJ��:TPcr��FDDT&�*a�ip�`���/[ʀ�K=���~$�¦P][.�~k�����+k�X��(��5ű\44�R���F��+������B�ai�0E����@dc���̦����203�R��o�9|f�Y���:p�{��L����c�����Q��0�L߿���\��	�	��`Ya�g���g/C����`�7����j
z�w�5��61�D#�f��@y؛�Hq�@�\�W1sI~A)��P(�î�֐����g��I��2��`Z�So�B,n���R�-���	8��`�$��f#�:��u�:3�6%\�ĳN�i��П�fDK0�]�T{ۤ����~�8'��� ��]H���e��n�S����	��$0���R(��F5^��a���Ӂt���>�7��y|�٠���hэ+W��`j��i
q���\�a�N�y{�e��
I	��φ����:���\�c�YL��INC��['�Ε�[܃S����������z�u�o�|x�	8惽_��?ry=��<�¯��g4)��{ұw���y]W+muq��͔.�D0�%ib:������wt�#r�	8}uAtf�t�����;Ӿ1������G	��R�6�X<D�ݥ~7=�
��������s���)x ��|���߅�䕮�҃�&�7.X���=�2V���/�P���
Y
����0��O/ì�0�]'v���6s|r�~Yf��ұ6��Њ���m��!���F�+[g�绩�֠�jl,��:��������$n#XU%@$�E ��4���>$�
�������|��RK�p�&rNK�_�P��
[��a�~��V�q'i�������{��l�LY���1�$�Ƭ�^�--=���l��xo'Q�����)Ѳ���d�ni"T;���`?���W{;�R��)�9"�q:�Z2���btM@@�W�+i`i�I�B�x_�#?5��ڼ��]Yi_� SQS���e�֍�b�y��ݴޗQ��$���b�:���Z7g���O'�}f�T�~j6�-�u�q�>�ݒO�A�>�{�_�1�n<�w]y��v[HUagWV=�DQ���i��^G�$�Ժ�7�c-s�t�+��I<)x��:���h��NC���:҂X ���H���%IB�Q�c��J�ϮS�Oi��F��;�A2� ø�8z#T�'>{6^SR9�ڥ�R�}�׻��֋)��xl{4�ƺ�^�'8�ߺ�=�*:�ྞ�|?v�C��/^I�=��nS�#�߬�J��0E!�,L\O�f�fGu��zfJ&P���E�11	NiS$�7w<�U�X3,j6f;�ISg���V2��{OzeO{m�`^�V!�e���(z�0����U��ٖ�T_4�ʹ��'��W깁W�s�p�oǬ�ꎶ���1ωLƻ
�
3��� W���]�8��"2�K���q�j�r��P����a����ci{����>NO7T�3,2t��l:�G.ֵ���7l����|E���餶��=ǁ���Q�5uw�z�]���&>3��nl0f<\@K]�,C���q�~��98�&v�3V��XA+�����ی��ߕd+��J�-}�W>?$�l$�����D�m�ե�W��uv*&�K�z�j�m#��R��tܫ�Zߖ~�j�&$F;���t�'�N����9�a�&!�m�(N�-J2jcp���oRY��M�F�y�4��&��%��Y1���Q�^�C�7m���������݆�_��ɮ�TJz���P��
�Mϑ��Tq�>�& P��,W k��_PK   �	DX	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   �DX��dI� �� /   images/aa7df784-6767-4817-a6e6-80fad30d0eaa.png�eTѶ.ڸww�nh4���4��-���@p�[p�4h�,@p{M�>�������c��FuwՒ���5����j�X�d�   KQAF �� P�a%vN�U`?_|u�=�̽h\ܜ�l�4>.P��� �쨱�����:&a����-��+�p 2k�P�����#����?64�>s%��*q�Gq4^�G���)�ө�
L��Z��u�n,��4Bef��cz��J�-�D��b��!x�'���Jm�گ]M|��|����99�H����zTXw-��zp'"�zdK w+l@F�j��/�VZZCQZ��؁1��,��E� B}NI��'�~R��,�2'Q��-{�/��Yq�٤�A�OH(AD_pM�	���n`G5��+�M�6ղ���<��%�
^�}R�Eg���"\��SL�**�7=H[}���������s�������ȴ�@��u�9�3Δ���^�����i�$���kϛx����x�A�[�c�.�Ζ�Vy�]*7���������wO@�Y]7�2JItez\��� a>-�}��Mj�{R���!����:
	����~��K�k��x�%�Ѵ`x6?8�|�'[�u)����>)�~,�MNv��j+���y�,V����,Պّ7���ظ{Y�8�B��i���E�:���ޯ����k�����-��b�fv��0��WU�8;r�[:[@��] χ����9��Ac��u�;i念�����S��HCml|ݠھj:_{��%�����0��#�Ü�����]�[��/]a��s17��&��t��4��nP0��)�m��C'�N#�fi%�%#�O�;Q:ann///./^.g7kn���7�����ւ�����ܛ�ɝ���?h�@�!n�.��N4����o<D��`�4�5?GU��&���O)����m���r;:r�kwYO��}w��rkAݝ߸A���P'�%a	���.o���c	�:@aM�a4@�6����ƿ������o/����������zn�5'��������e$,�y�<=EQ���-�!���/yyx�ͭ�8A`^N����X�i�o	��@x���������L
V�e�#ᱰ�
	p
B̭8�@s~!NsA ؊��JP�_H���¬���_g�L�F�F��,�) �r���9͡�|�<����`s+���,!�r�n��0u�:�[C�]���V<\XRCQ����?%�V�0�u�t�r��*[G�����<A@ ��		���i�us���3U����oͳb�ف1a���_|
K�A�=��t��D�I�<���jU�CY�{�˘{@aD�<`a �0�	��A����������������Ј�C�
���}��ç������ǭ��?nh����9�,��{B-���
bc�d���/��_���� �/�� L�<V�B@A�1�ZB,�,`���Tܝ�<��ݠ��09�d�ʿ��a���X������B��p������,��r+�����?�K�y�\��]�H��ߡ���?|�g���A�3��� ����A��LA�`�*M;�W�`�����_���n����(� ��8@V	��CQU�'<" 	�� �  �(�H�x/v�uC�;қ��^���(�P+�*af)u|��$����G`��tTE��M�C���G����e�"�e%V:�*��(B<tt�`㫵k����C~'��/_Ң2D���ge���ͻ�{[ߣ-���ʀ�����mt��k�<A���7�n�!�z���-�S��V���\� Ƕm���u�';;��ǘ���}��Qa� ةdN��R����'1��p~��ӄ��޸�9�"OO]UTT�,,��:�x��d��0�]�4�׀a�w{5���w9As|g�8MD�k	���p���-�2�#�&�����ݯɪ��5D~�,s{2 :ӣ^~�{s�������
be��wy�;>�y���=}p���2�I��4�VbE��{���Z����R4贡�����-#e���Y\h�C�	B�ʀ&_4#����H�6@4�Jl������%Y��;)� �@�}���K�R�j����%Uȋ��m10-�V�i2�8.�nz �ֻ(E/I����s�a����yuw}��k��d���0>~	z�"�l�K;��@�d����/���(�G!	J�R��*qp�QՄD�$X�/����T���*�ѐBt(�2�ۏ3ߟ-��lӴ���mpp��o�T<nٮ���qe�6���`~����`�b2�olX�If�K��/\YƕfǕ6�P�����b=���{�D� ��[����Pd��R=R�׉�{h	1�b(����plY�^@�&su&��+�@�5YZ�0���VC�h��	%!��M�$*Z�K�9b��(MZ��ѝ}5MI(�P8ΰ;-b�0��x��H��~�2QѼ���G�AR�g[�if��d���%��ܻu���ge`�\��Q��� vw����E/�a���[��z�H<��֌<���?�z��P��F�`��t��|��q)A4PN�����=��~�5 �z��m���iD�wP���� @��Q2w���s���d	/�;��7��u�Z�V��(O�~^��ÕS��V �#/~�|{��������)t�:�b����"I
���R��IO��`�r|�0�@�(��c� 	�k�<thZ���B�U�䒯�Â�G��J۵��!J 3?�fR���}��뭛� ��]�@䏺�Y'd� ��O�E�S�H�r��^:��.vqQDy����'�y�3���O�v���l��323]m�Pi��<��K�cAv�E\�k��q�������C�H���?P��H���1���Ce��f��Y�0�r�Ѫ��ZR�,0V�-�i}�*�ۤ$�@�����a�x���U��L!�E�d)�����/Vs��-w��u�sL"����Vw�f��У��0�+��y��x9�T-�/26��d9��X��#	,i��S���&�2 g���LU����x�d`X^6n�aӂW�p���V��Y��&JطQ�l��1�Em�P]'�O-�����fEYn��X��|M W��ΈoU���q"��N�J��@�E�o�,R'�w�\������^�8�u^���9��;�u�b���9�~
�ᓠ�1�c���ĘXu�i�&kFi���Ve� H���=ۭX0ᬬ�J�lSUy��t��De���t�7�e��C��Y�fsEE���"ɴK�~�ӿ�z|y���k�C���_�x6�*�N2�<��-b�|�+��b����N���gW[�I���tƬ.v�z�݋�����֚�ɀW�9埻 aJ���B.!H��dj��@��b�zt���BB%�Y�!���	�:�R�"��R����4�����Nqy�O�ļ�&��r��C
�aQ�(!S�9 ����SO�S�����5&�0�'�ycVپ" ��2�C�a�9�W�H�)�b�����ȩi���s]������$j�Z��)�����7b����8д�d?+𵚫"
P.[#'�+����;Ts[4$��^"���YV�B;���(�S��!�����Dgi�.O�J1&<tZ���F�3e^̟)4Z� y��mFn���@���&��� N`a������f�s�q7�ܩ���j(�KO3�B���o�d�-ܠG,���𧔑�o)�F�&M晣�Y=7� �,�@Df��Bhڼ�<�}x�6>Zة�������I3~�I3�$+dE{�X��Y�����#��b;,e��%=$�1�7[ó�9��I�\�3E�n9�k���
t��{��"G���A{Ϊ�`�//Q�ɝ;f����Y������B{����Ŷd�b�[L����p6�q!��G����b�Wk�+C!/�P]h9�l�;�?g�5�g���%�I��h�^A��O��Ҩŕ�B������}�����N���"���M	*���,��9�,.���)0�(W��B�Y�v��!*�u�	H"��6I�����i�^':���d��P`���V>��Di�/L���pH���r�wG��a�7��]�F�<l��B֘1|�kJ8ԃ��@ˠ��k�`��͏�DW"��v_!<�3V�쟀�ځ_�H_∶c���)�`*f�c��%ef�Q4�Łh���+?��J���X_��DJF����X�X�+��IB���%�V̧rE3�<g�=j���r��������Ѭ�~x����>����MV�
��#�V�!M2l�k��\���	��8*o ���L��|V� ,��8�K�-�[|KK��H�@�SB�r���n�[�B�h�I+�����a= �Ȧ^߯��B/�m'<?��i�ճ�f(od�D[��SÌ;�?~?��Gb�D�Ϫ��u�'�w�x a �6EN|\yI;��<�9��ؚ���l�����|���]}��̫�,E���`�K��n��s �~��N��`�0�%ℇp� ������ٕ߭�󌦒�>]���/6���*�ڢ�T*�5�@	�$�ԇ~�iR{Z��sR*yF�_�v1A�$�B��R�����i�3�h{^��}`�ό�|-l�����*+���@.VM���ZRl�͎�5/ce���K�s��.o�b�?�m[]Zgn/�a���V�b%��0����H�~=x v�:��V��6��k��و��dᶰ���%�������hZ���B5A�͆���8*��B���*9�rX,X0=cG)�����A�(z����0AEڧ��;k���4[wnB��������Q98K��/��������YR%��
�g܄��|�j��F8����ӸfA�!j;7�`Ul����-������ص�*���rݎ�f�x�&~V�*`+���Ŷ7[�F�OK��r�WI 0�1�Z�s�UF��.'Yo/�^V��/>|�)13�7ʗh�-�jR؈	L���(D[��Iл̉Y��k8Q��P�*�+P���Rb�:z�U�No�.����F��t��Q6���*8*c�f@�9�+
�ݮf��g�(��ec?]Km�Ib�*��l�@�����h���	����թ���y�5�P����Jr�0Q���]��\{��w'�j]�#O�w� C��Q�@�������~!�������D�R�[��<�7�L���Ɋ�B$�WS퓁J�#�B�b��qÑe��Ur�bH��"�4+G�%J��������t_>�(�WJ�ʝƵ�I�O��2��@���z���j+�Z�P�j�؋��k�F~r�/�б�g�yc�A�j�Ok�H�Oy���2��;�j�=�b�+=��H�q��84[�\��7���̾ ��yDf��ǬR��a���7k��t��%�>�ٖ�{���7�a8����O��{�_.��a��4.m�,p�DzW���ޱQ&�%��O��
_�7��<����Vqk~�s����q���h�<0�ES��U˥׳���z���}�w����zP{F4����C���M������V_wKQH��Py��s�v��������h����8[>���q~|o�@JA�ɤ� �	��k��u�Y2N�k��o|'�=o�O�!O�b�zw�"�q�Q����`d�L���w/ݍ@�zoH�[~ŀ������&�&(/K�
�K<S@6��Qf]!ˇ���+5�T��5נ�ocMY�Huk>���#O�;�)}��"�3��}w������.��g	����e۫�S�&�v��A�_���F�*���<ߓ��������x�I�ӝ���{4<�.���*3IZD����t�3N��b���O�2��X���?���W.=w�[k�7VFbZ=(���w�yĤXy�m
�|Qi�,;�h�:%t�i��Ξ{�l���hy�i�����S;z�o���e���<�I��K�ė�?��JQs!�>�8!��t6���ܑw�Б�����`�.�Ѩ�l�꽲�iz��z)(�ٱ����޳^9�Ǉ�.뾟��`~j��������S�ƕ#�:T�$eR�q%����P&ga��M�V�j�a����Ÿ�����(v�����Y�ɛL9>�Q��²/�<]�8h2xJ�le��Z�ؖ�nm�X~p�R��5r�REY��Qޭ��XE^�H����������Ȅ���6/W�Z'�Xneţ�~�w�c�&�B�.� ��R�k��-X�k.*0O��vM���-���c?���/`�a��Wc������gZ˃W<6%t�\�J٩v�mU�}�[~R��%��w
_�#ǫm������J(R5]��Ȯ֨tD����Z��Oei�G��]ͤz�*��e��9r��M�;5�+�$8�����)$$+˛���2P7z�_&�jVi�yO�'�Ͳ�4�Q��x��Ӵ��DZ�K=V5tqk��G/�B�� 0��h���z��-����s��4�Q3N�
2�$�����7�S0,F�nGGG�VR�R��!H�XF�Dk�IT���sŔ�����TגI9^q��=(Eܒw��M�zIHx٦d���ԋ�W�V3s&��URE( >��t��+K�Ά��}W���$:�&a���t�-^���eG�Q��|AC~���w1���n㧇kTE6�"��;���$Z�KC�y��w! 4y�l{���'O�(�p�`3�:�^U��}�}do{ձ'*�����xM�e�����cH,�)�E�Z�	�uW}�����]�,``���W��άt�S�Ш�c�\���)�q�44���l�"N�Ϳh|ી?F���@d3?<�I7ץ�6&ܚ�r1���u��/�Gp�[��Ku��臐�g`�t�'�2��K/�����hO����|X�i�&W��JdjN
��k1��V]W��ʩ��|;W��<�8
�ksc�ׯ�ǫ�"S��K�ۇS��&Q{�'>X(<h���RX�:��^�~0r����wG�R"����]S����������6B�XCiy9����w����7�:V֗#>�O���Hb�Тzt�-�g��L+�F������z���\9�����O|8P����/ieJ_����������������� r��8W^�#z�[ ��+S|�����*�f�n���%`�U1�����0�P�����)�.k>{���TB �h�&��7X�|�Ga�;t$AS~k{��7�LLL���Să����xs ��ո��a�D��s@��f�2��,��+�׈C�d��T����o��ЕX�ߥ]��纸L*�׳��_�x�u�����/��G�HF,�;>-��B��ֵ�.��o[%,>)؋��A�Tu؁q�</n�J��\gĬ�|�*�jJ\�+Z����d�	���̔�Τ�_Zs���+��$�˅�3G��]R�J��p���B���m�}a�о1�.�=�b�ۜ2�����=޻�*f=h��B���"��~.m*���9��qN%�7�n=��(Nrt�L��#[��b��՚��1tuo��!=ӟW��盗o���b2��Z4���r�4��x�߭�4Wmx����;*��Կ|\sw�V��݃LW���#y�
�{j�h��ɱ� �S���"�N�Җ�l�!���9��F��	���� v�7>Q��鳈����7�UK*.�&��[�"ܙ�����퓄����iמһ���zf�^�7�h�0�)E���1��[E�(��]����-�d��V�ϗ<�N~��t#�U��=���vX�Ǥ��G�R�1��mm�������*�Mw��%�%���+��Y�^��.r��+�s�̩�OPV脔�r�Gt(�}���vY�*�*	�C�h9뽬
�����(_�UT����i�$����'M�!)�<:g�y�_�-������J��B��[����)����/�G��r�m@)h��k��49���ߡ�()Kd~s�C��x>�|Ӫ #/�?Z>\��^O�u(�V�V�.V������#�L ��иw觲w$*�S�"v�q�Y��[��YѴ`���Nt�9~��R�ՙ�`��!d
��/[���v��w�W�����
&E��0ܼ�^�1�����y�nz	/K`������������k��i�fس�,�뫾�=�K�*v��ULA~�H||.d}]b�5��y�к�#w���D�s�3����~fXj	qp����K�)�� �W�x/m��C�l蛙�jP䋝���Σ�����1A�YWҔ<i�����߈�Y���J�3���p�B�[�q�E��>͠���y0�Մڝkdq����H��ej�>J�cR��e���G���b���g���~Z	�-&��N5�II׆��?��F�z� � ���J[����͌�P���ʳ^p~82�~��.�c,Ɋ4t}Z$>x8�9)��X�'�a���<`Y؋��>;.F�b$���u����d*WT�qN�ݢuԾ����$\'}�wb�!G>~��)WknLr-f�H `���L�Zbb"� Ѝ��2(F�~��6��l+�cقSS#h�<�0Hg�֥�KN!=,q ��H�}&���=jߨo���s�����Y	'��٦��ce�h[6���(���izeGu����d��mT�V�f�(���=����W9���l��
�J�e�J�k>����լ��i�%3���`"/�BP�f�L�:�)��"�/�%缠v�`.D�T�
���A�ϫ��A�R�~�uҕ-��#��=�:2�y��W��d�:�t��\�]fV���T&,���b� I	c�f���N���xi�໛5&�
�T�����4	9��U�'+<2UE��o�+6�U���ǻ�"�����#��Rc%�!ӧx�ux{qu��oQh��xT��Z�q����쌩���k��Q���Z�h�
�l
+
����_m:��;���O���r.���|��}j�
ڼ�{��U��0�Ź���jD΄�A����&v�������b ���(�IICCnTa~��a��b� ����gF7��xZ
��h�cU<��9��Aqm�-cJ�*9��9!x��m��7Iŝ\�*��V%��4E�"�Cl,�I��q���e��+DUB�Y4V�b�ٚ�e��
�K��\+�M��ks�B�i��Z��ppZ%�?�(b�w�Lq�O �s��Q!��0E��6$^�N�zR3�~��칛���o������V~�%����o��q�O�`�%.1��/lZp鋲���v����I�0������6�9�ǹ���SmS�< �ZH������ڢz���߶,�&" e/_�W��,�)���	�س��!����I���;A�;�!M㊥'����˄Z��(���lS�6L�L�`7�f����Զ$h�n�(�w����a�I��چ?��q:�#�J��h2N$ �,���~P�X������}O��~X��2}Tm��|�6���` (Z�τf8O��gNm�|���u;
����Hc|+�J��)�;��Tu/�?܅����J��M/77/�����2��!��bP�Dz:��mGk�HPbS��Z]����f;?$2=,1@U��k�tG��3��q��{��.��:F��Q`i��=ZDE��I�x������}P ���5j>�����V��# �-���b���H8K��O���,�=O.��xe2�Na)I�$�Oʚ-���Bu�}�<(�،��b���CC�Y9a^�w���q:6�_LvJD��i�Y���O���9��_�,�]7V�>wz���q��1*����D?�������+ePU��8�3>��~N�g���z��eY�C�H���J?�MGI�a��H"-J[�g�	�:f�OD��{����V���U�ȝ֗|�X��J������mg�pn���la�����U��x Pz�j�r��,IVB;'�Z ,��P-�8�l-�d�5�mJ	�Q�K+]x�;꾾M���"�kS)%tEBT��f�
������9P��f�Ɔ���C�C�e9��F�7�M�W��;��L��}����%�ٺo�-��i����~ʋW��~���q!;���H7��  �g��^���]V`^�G�y���x@C����H��B.�B=fN��>0�w*{*cH	��	�Q�6=.��?��A�����Y���+x{��쪩΃�&׮&�����2/rKNR�=���V��ux>���p�Nj���8d'$�hą|	�}A�(�>�^SWZ���!�C6wo�>�T���� �c��%ݐ9X�^�5y�u��.M]�j�}�y�"K9�1s���=h�9��f�o�Ь�)�<J�إ|�C�v������s�2]���5��>:��=�<�֜�+v,�T�LO��J߯�b٪u8Df:Q*���d[tey9���sN��~�����?}B����%Y���	+x��y�K�c��_��֐�@N�1��ث������c�N` !��\8���C��~T�{�"��B �vЈ�JZZ5y�L�"j�.��EI�hps��M8��x��vF���?��4^�*fEhh�1?�����9n��SK��[�n�'���iq��4�'쫁��a��]/Մv��Q	�9r��0�n�6�k����w�l���������_���x�$W����
�TQݓ1*B������| ���V}�-br���Ō+��a��SW�-�eAe����>�m�>�NI�j���X�REs#1}�����d�E6C�$2c��%eǉ�IB�T���4-����f�n�SG#�ς4U��J�e��Y%/�;xkQ���㍻$:�69:J?m�b�<1�E��j9E����i���J��&��$ �||0���פ�
k��r5�����FE���"�Li����!ߛǫ�u�}e�>�Q�z�Z4��SHw�O#���
Y��n͗�+%�|���s��c!+���"�����6�(r���@k���sH %GH���̐YZVZlN�k��	�ָ�2�Jû J`���u���L�R���&];��	<
��j�b?I�E���T@1����&��`B�i25�գ3v.����VbA(�T��Q�$�q>D�����������ۧ��'懾���Rgu8�O��w�MVX<S2���m�����o�h�{�MN�U��!0��HV�B�]TФ���|�{a�Ǧ�WA^��	7ҽ��}��(��#�I��������e�E��ۦX+f�.�?J��F���M���]x��)w�%n`����"g��M� �?+2�h��\JZD3��Lr�7��d� AEyK�j�}56�h8�{�3lQ%k4QL�F�I��1[���?a�xI
	55
3��&Ok�˕/B{9a�\m�{���C�Kn;�;��K�P�����L®V�[��b]�T6��|^��?x�ON"�;o!x��źɺaȽ+h���զ���f	���&�4K����Ґ���@5����F�אN�ђ� =DlL����0�*��f5�#}{M)������HO ���WdX\:B�CK�8�2(eY�Bf��9]Ϗc����A�r$܅Ղ�8=���<��ؠ�Ȧ"?��Ma��88F�,�bŘ��a�1�,����7`�m���g��ż�z�q��|�&iӼ;��bF?��Sl"��H�<��z��r��j��j-v�; ��Al�{��j��s�VN���k�^	Rj\ ɺ®�EN>̇��C?0����*V��e��rD|��:�r���\���GS*aQE��L$��^/��G�����z���4�}�L���/G(~[u�iR��EZ�b���;F�ʗYS�ڕ�hY��_ޫJN�I�qP:A͙�	V�7��t/k�HL��O�sz��5^���&Xe	�>����$��1ҔUTO��&1|��z �	�7�� {O*�OFSTqt�=7�^��M�"gP�/��'���Q|�J� ��6���{��d-�PE�43c���+�/mL��h٩��s�#�����]H���6�Ҋ�#�:8�����}5ij�`���-�����i�`z�_#�I:��Y]@|���jon��A"�7ɞ»bDpxVRe�'ۆ���Uj��%�ZkR�=9T8VY�]p�@
J�W\��P�#�|�*ϓ���E�7�G~�r�n�>���h�����x�������r���[�+�?w��l�^�[!��/�F��Cu��QÓ>7��L�p��q��3?
OJʗc���;�6)o�[���2	�9�����ز����텍�˩˴��Q=�_�E>��ډ��0�R�s�o�Ҹ�&3Pd1���
92E�~:��(&�`��88�iT����5��������ލ�Sp���o���B��r䌹�U�qR���H����C�-?���1���v�Qh���VO�j������G��;'p���U�����p�R>�{�#�'��FYң_�p��d����n��^�0������@�{}�_߭b,I{x�'��M�r��Cd�!�O㋚��ȵl_�-<~�e���of�ȵ3��l;�r�	���<��:�6v/�9�s��5�H�i���������dr�
�T�c)��0�7��$�,PX�q��� ������nj��!�y1�5�K�����9�
�g���د����z�l�)���r��l��畟^~���Rc������K�[��XP�qm�9+�Տ4�D�>m�r�d�]�&�.n���'q��譐��,��y�d6^L���'��&�3���W�[=]p&�w���n���21]�[��Oqz�
s�U!rE�3�a3|����t���o���D|���V4���(�G�G���cȌE$q�	j*����N(e1�@���1�Ȼv�v��"T��Iӛs�m��ox�'�&�`q�{��z����W|����Du��Q��X�� %��n�e%T�/�HL�7�Wx�)��LF�Ԫy�%��7�~I�f�W�%n�و�B��bY�����7�?�B�6�j�6H4�@>�@+6��}>�����;���AQ��̯�����Ʒ�}�03�s�X�8i���]' �*�V�L-}"4NO����L��x�0��/���e��D����}R����J�~���١T#$9\k@Q~��3�x�xI��r� WE�0��0���)��5��/7�Qsl��Q-@ ��Q��BV���bQ�(�K�*A�m��t�j^��@&����̘����ԟG�W�X��"����s@㞢d�mź����!<jHh$fO�:'}��j�t�GB=�x2B#�~�?R��� �D�3ꖣ�'�S��5p��,�|�;{����!�9�/<5c�s�W#���p2�Sr���������2���;X��0�s���srl�하(�k�'��V��~LN.�(5�W�Dkx���"�pp��.ʔ5:m�Z5����}�9�fDIU�Da\�L���04�B�5
.,)�8�����3��I}�����k�~��+	��3 	���CS/��o�}�>�ښZ��ٝY�7<�RK�hݟ)�P��,v��֣U�/Ve��`�bҠW�4����i�^q@�e�-$&�,�':i��}�F�m���1�  x4��V���RތOB���~�&�p���ֿh����,�H�:k�����.+av��%͚`��͠6)���,0�iU��͉�x2>����x��-�G��>�6 w6ϋf���y���cb��1i�.�5������Ǯ����l	�V}("���W.{<�$��/jX~ݜ�]z�"1��%�Y�N��P�~T@��7΍������'_?�T]sb V�r��A�Gw*l�
E̼q��u>�rq��
���r�O��)�h�F��gJ`�S�re]�A���ͥ�%��81���?<X��E6m���m��`)�6Lw��5B(����wlK|o���U�}�Kڻ�I��~��w�S\��Is}<��)����z��1�\^]�?~�n���� ��� �XR�'ε+�Mx��19�`-��^c,߱J8�������Պ����H�(b`��"_�<<m��4|�,�s��A&�q�=�����Ka��#���p��n��pS�3�$��Hc��5T��(�c������t�ĦD�)6�����nc�M?�����ǎ�~I�e��w�[䫲\��J\�!��]�冡����i�{���O��\�������W?�da;���,r�v&�tкʮ$,��֝]��s���	����}�����)��7����Q엊��%�5�=k�E��C <R�6��š��C�-^k@�ˮ��}����u��' �ZA��:s�U-#�m��{�����!�[zS";��wkO��gڲ��e���埦(8i��%��h�P?�Rt��;��ۙ�� �m��p-�P�r�`����PI�%�xݔ��\�/�Z���K��GX�C�����N�3�n
N*����N�'5洗y�1�cea��üʥo2�--�D^�X��R�#��0*N�3��n�����H�H�Ny�?x��FVپ��"���xɋ��DF��ϗ?t7}�C5+r���"JIR�	+���[��F��ԩ��{q�&��.�<i�amp�}�U�z�<5��U��@-�z�~�ʹs/��#*W���hJ.�`L4���.�u��?�����(慟��݀�/Jk/�5�G��_fx�L�g��0(����2� ����'��U��غC�C��؏��؛�@�@ꆆ��W�?��H0�P��[�&�YJ�wL�7ܑH�4$����}D%1.�
���b\��$��+ɳ6�Sg��]�Ý������DkK[�y�f��W8�ɱPt'V���E�%��=YKhhl,I�?�?�о���r��F���}as�L�Q�������C���~5OD��9l��v������� 0���/��@��ӽM0i)���TOQ�� R��0&Y1�̡
�xE���ڵ�X�X�*eӦ��&�	������i���|�vSE�H���(��P�Y�/B�Q�6�˱��ͧ�G�U�ّ
�� f�h��0��P7g�°�8�gxK�	U 0I�,�Tjr\uzI\JZl�g֭ҏ�N��Z󣞜5���v�P��?JF�9e\��Ai�_�4�*�=<:-�{+��g;����h��D�7t�ѝrZsLŔ����Q�F��W4چ!Z1��*�o�:M�?_[t_�,Z��5�L8���j-�;L�EOj~D�B��rjt�����D�	�۾= �jkL�M�Hяٚ(���b7%G��~aӨ��L����Ϗ�a��Ӳ���{P���Q]�rgH����M�a/
�����#�q��9����Ư��/v��H�����$�̲�;j��h��pl�Ԝ����6��M.! z�~����e�a<�w���ٱ�X�s�+�׸����C�rbRt�7t5B��s�A��A�����qxCoi=�����8	�Rq����lՌT�� Y��|��`2�`��J�6�*ä�Y�� ����D�Naq�n�`쒝cH�6�0�� ���w�s ~���#s�!O���*��q���[ԃ�B���������  ��m�#>DLώ�dй�DXv��C�ܹQ�욧���V�^�?��hZ�e��1Gz�s'WG�
Fu��]���Sa؞���OQ>9*hU�̀���,k�����N��X�We����$�VG�H5��}�9���2�q��<���fT���I5>��PwA��'���Mb&�Q��,�<�4}`K�%aP��R����D���J�$�SwP&������[VX�Y�kJ�#߰��J��V�G�b#��h@����m���/_�@���s'��
��?'j�AuR�%�K��Lm�-�Cp?�y��d(�����z�-�ف�HsG�wך0���zbv�N㍜|�.:DM�N��i;D%�9L�a��~^�Л�*&�Ы�;�7K�#]�������Q�ɡ�6��%��{q��畦.�����C����ה��Ȳ�DjJ'���|S�_�p8���m�٭S���D��� ����<<�N��	�7��iv��p��d ��`z�#iO��yk��U�ӫ����f\UL0q���� l���4.���Z�	���=����M��0k �)�=Sg>DB2'5���?�Μ \�+�(����4(��y�.��"\æ����&o�gZ�L*�7>�p��#�R�	��n���Ql�/o����(�7��KO���j;���<�f����f�v���{���Jyt�J�- ���r���ۨ�`��88�i����o`R$?^D2�A	x�|��p 0+?y�V5��Iʳ����V��[��W������$��RRa�֤L�L����G���+>~��q ���wM��QK�!R��.�"�2�[ky�8�� Z�)"��O��!@�5i�����1,��f�MU��k�+��Y&e�����8ϗ05C�EV��}�ZM6��{Ub?J���</��,Ph����Z,�����<��Բ�d]��P��A'C`��������N]7VO�iO����2*��Y>���@�ஃ���	�n	���Cp	�!8�ww�o�����s�tU���[\i�1�9�%}�P$�[QY��yPQ�ހ:�_PX QГ��������M�dT��;�pG�>�x/&�@*�(Q�2��ئ&@g�/��[+��j�S��Ce|�MΠ��K����'�-A�/cJڋRO����Q�B+��R��	6�������Q�-��10�a+	F+����{���x��*=pp��z���4��Dm[cѬ�Ž��	��P>�76����2ή��
!*h��YH��0s������)�c:�+}�����~�毆���f�������e�Bhdڲ���݄N)hث�Ő�N���?}�Hը�RMZ	h�A�D�H��0��x�lq��x����ь��؜��yHΓ�M���¬��dZ��K��]�{`"b�G#4JX3��v��9SB���-@�T0�B�Ā%I��]S�5����,�x�\ݲLv���~��W�b$���������`����%c��T��7�W��O"ؾl���:�]�~+��r�R撟�y�'`��*p�8\ĺqY3y\�Sw�xD����n83�W���q�>�[r�^�84O��p��@��_��N6�_�w�m��q*�I�X�纷�ԇ���ZȏU��)1l��#$��i�o�[��y���X�-�cT1�[��B���ngȯ�ѽAg�γ�硁q�{�}��n�4pV7ܗG"|EV}����Ϗ䙗vI�?X'+˧� Ӫ�d�r ��nD0���9ؐ�ɶl�kC��t�9῍kfSn\qR�_bm�C=\�`s����=��S�s-�4A��������� ^��M��#��jX �?W�q����C��\5u��9�2�Em��N�he�	���2�-ee
H-,K�$Y�Z���?���X�Հ#$�7�iKH$7���8��P�A���?]���PӨ��%��F�J��s+⶛��fZ̷W�1���s���v�O��g�/�m 9T1�#���J���}�-3]"D��b}��(}�G�z!�8^�^FE����۬� ��<G��	��Z�N!�yu��}o�8P�v��Z�����7�ci9��sΥ=)��VV��a��-�T�񯷨�i`�2N�����K6S�"Ϋ}���0t=����PH���ԥ��J7K�e��C&_���T�	��*�T�9�9�`Q\=0�A�vB��,�FB� �k!�--�m2��MV����j�D%�u��\{��|���TcF�oM2�	)N#^���JP������7�ri���uMv1Tuu��)b#zT	P�WmcU��}�PdS)d�9W4k���s&4���ҫ��=����l�P%7GbNM�b��;(�*`Y4l^�Jn]i��]ͥ���fW6~�"�5��q���p\<�{��r�Q�Jp"L�G
�o�tZ�L���~BŰӁ4�-/��C��2��bS���$F�ޖ��H�I�4%Ʋkv'�,B&-M�ܑhZ1�ۼ-KJϫ�����Wy���;h{"P������_k�3ě)�O�����#�S�L:��y�ua��XU��]:�	>y��8qY�E���X2����V����4\:��:�eۻN�D�ɤ����Ô�a��a����A�$�� ��)Ș��T�¨tJ-�ˇIK<�E�GJ�������Ҟ�������S��+����d*�iZ9e��:H�A�
�bW;q����rm���7	P�y���g��]d�p��RnR��;� gc)��0�)90�,�[�/X�ai��x$1Ѵ�����젤�>G�"A�}�M3�
��E��4�ܓ��K�C�n�O3���,�-���v[e� ?4x�~��b�3��R!
*YrLi�����f�l� �,Y"g�W5ȅ�	a�s�U���a=,>�i��ՙe�D��ڴا%.��e�i�d�@5��p�q�bb.:��P3��@��ATJ���D���Bd`Jҵ���9�|[��N|��c�j��%��l�e���rBUP�:�#3�C������!�6w��г� �T_�*�G�^(T6�;/��L�1\���G1j?'w^Ž��|pϪ�=��W����6;�xLx�]�(dq���F����pe�dy���:�N�j%�ǱP�ގR席n!�:�K�K��3o�a[0c�?c�\�}K�����Z��z�Xn{��1��6���}�'�-wܕؽ{��/��tI/x�w�6��L�������$UuT�Q���MP����Li�V�9?��:;�����,��n;do����_\���7C8�"k@���.���+��sK	�o��l ���	� %獟��k�ZU�����od W��wN (��y����w�+3�#�/#�!H� ����,]�\"'Rs���A���h_��_���o�	H3���+))���
�����Š��d����(\���Q̥�'{�=c�"��,RpHd�d��3W���u�ƽ�]|�F�z�'�ئ�B1��'���Bkǃ��?�
�3�"�PIf&�-�����]��բa��i��J�0D'a����ŵ�B�a���C�'��
�JQ�T�=>� +XJ�����n��f��o��a�xZ?�"v��$��Wm/::�#>��t�e���ЁJ|��ݠl�o��V��a[��	�ϔ!>�Ka�c�!X ���E��� :X0��5W���9����z�4�c4�y�6���clƵ�G(N2ߣ�u��3����It��y��!0������XͯE8(�L�\���+x��U��ڭ��E���$�26�BB�1C�ގ��`<Jw���7(�_�UF���ߏZ8�c��Nd#���/��F{���K��3
�O[;���PC�RE �G�;I����#�]��_Q�7�|�8H��߱	�1�=Y+����O%;A�B)�h��؝���"���'��i(��Xz5Z�囿�ˣ�R�W� �X1��0�	IM����
ba�:2������M*����:��AdW�<F�P�g�߻��O�9������P�@~q��Vu�Z��5�H'�&R�_Bb�@7T] �}~=k�<:�����i���{�W���br�]][�w�V"v,�w�!�<cF&�p�%c�:����ke.���Xs��w��7x,\��J�S��d|�,�9��MɊ�p�f��2`(������=>�c�f�Ԟ��y2�k[�l�P��,�BblA��K�QLʅ��|2"Q��$v�w&��`��O�a�{0������e&0���+���K%@��N���M,�2)�ho]]g�P`5<�%؞���ˀ��>w�g���"����4���`��<��,8�DG���"c8v��-ȶ�����&��C�-���=X�;���]���+�BV-&666�x�	 ��M,�2.O��0D�����VTn�%��Dpy}�����'�����ѳ����q�~���f�۬lzzzw��/tw���Wwe��6&�d+�="�Pf�Z�،�5���졩�}��c���t3ξ�o2���E�����;��%�ǮA_�G%�3�t%��b�����[k_#����;�4C������(�?�X�=�B�K�g�jFH0�8���1�oY�[��Kcc=7Ph���I�>�K|���鸐�<v
$633�I�]sl�,���<�$[�qR������F!���� �ƺAw�A@��P;)���=��#�w�X��Jz}���
�5,!��2��]|�Qlb�I�1��d�0��H<���%����9��t�#�feɺrq$���x�6 '�u�J��m󌛐�z���Ӗ����S2Q,��1���k�w֔�н�������Ωm��G� ��S���i����L�����چ�iK�0������Pz�	�w��*�]D^30?^����I
{�B�*P� N���N`�g~��@��[�X-��Xn��P�M�J)h֖[��wʕ��t��B�Ԏ#���!��X�RK8[�l��:�%գ�V켇�ҳ���ۼ��]մ`�3�����,���=q���Xb�Q�Ұ+��/��2�	�vY�9�mU����Ԓq��*An���:��f��<2M�����|{�w�8b�:����#������� �Hn���`2�UR���qקqʵv�����ϻV���2���+�D4J# oRBE�LY�̺O��6�w/��d�Xi�G}+R��U˴o�ĹIYT�erqݹ��*���5��U�x�Y��z��i뚶.�a�0�$iWZw��lSlN�̕��Ó� �r
>�s����+7To5��@Ӵ����;���f�8.����!'ͼy�ql-�c� ����J���*`�P�0d�A��M@`{����#�y�(�<��y34�Ų'�J�R Z6�r��Pഃ���^�A�B^����u����� �R�Iz�)���y~�^x���U8˄Y�	�4���)��X�E��9n�c�*5S����^]A3d�)���V�s�k;��~\i|���.�Z�5R�e�=��i��X?]}���A4Ů� >V�oP9cj��Tԛ�D!���,�&�6"n�r�<���>9�y�R��gk5�ˋ%-d	���T�����S����fNv���6�"F��}2��$��X:׹(�o�&�ط��qv�ڛÙ�ĀI��Ј��/Ě�mH��So#���j�D�
d��4۟_?^�
T��2i�7�L��h�oH(��`(�J��-�Z�(��'��[�D�_�E��= �N��ɉ	!��bA����uj>�tO=�wU\��ur�?qC8q�=Q��l>P_�w8=��~�G�0��<S!2O�P��s7�Ya�%L�~7��Y��-�hD[����0�����|ټ �dg"+Ҷ�V�.L3Al�OY�F�����~�?U�?>ժO�d���$?(�!7���>a[�E�8Ė6,��b��W��D�t�8�h{e��߬��T�Y��L�Q�I���z,���?��,v��&8���
t�]O�t������~��U�����K�@-��?ŷ!YM�*��26���#x���V�0��˲�qh����y����F.�ӗ̂?%E�8�Xf'�ks~��rY��}�B�3����o���N~���B��
?
"��N�?j!#���&��lW1W���ID ����2�j������B&��B7?��$0a͢�H_dia9��l�����u�"�-�K��E?�P��C���)��h�B�D]ʬ!�Jث��)�c�E!�����3�Z["���w��"q���C�
�b�6⪸z�ձܔ(�ݭ��	r����d��hK~,�"�y�Vlg��-�G��m�T�dβ����J�Je�iE�+-Əd,݄��ń����f�;Gq_�)�rtf{�Ǘ|�<���+��l�g��3���F���
��YGEA�׶>��+�l
���+>��	�C�ݬ����V�� ,�FK��_Q�=sz�q�}m���zu{��'�#yO���)��/(�K7�J�tT���V�=
�t�#YcTyc�iSTYc��X��5KT�M���@������[(��|�n��od�$�~d�,��0�b m���!�b�Y�Ջl|6! ���=c4뀨'H���O�R1T�i"�y��|��j���1��i��Q�.�,��o����>WaL�^ZZ::�u(o<�K�K؎��&k��e_҇ʰ�'����7��c.�<c���X��pӝn�)�X�=��`V��r��25���gӼ2u�MȀ���7�]����eW)�ǘ���#���e��[!�K����T�t��q�����F��e��RC�X����B���o���|���W]�����*�X���N����x�� y�P?�x{:�b� ��\���\q�~ty�k�ildCR1�������CXLR@��������'�Om�-SĨwb77��d}�%q�5�?�ķ�±�'[����yPǪC���p2��)�9u�j��R
q���nnn�4+M.w��NO�*�\�J�d� �x�3� �y��F>��	�!:�i��!2�@Y(J�0��/��kx�S0�p;p��3��R�,�r�b�6Gc:�}�,\��y9QQRy{����+�Z"����~Pa�cIl�ak��?�3��E�����mG��u�}ĉ���"v�P&�a!uD �|.��)�D�\��3DDe���1��B2vCx.��z7��O %�4���8T#�*9
����`���`|NR�o�r��}���%��� ���U�E�	;��ϭ�S���E8@��x(��|Ւ|�fTO�mx�A?G
+��Q0���'{`����<��B��n��x��c���� XNx���̶��?��� |��1��~Lld��'��X.�-34��S�+Ь̰T��rXi�~� a����P�"���2��wS ��7 �?�yk���͍��	�?�2
���R��b���m�Rs�1���R��J4�^�Z���3lO�z�b1�4T����:~%V�/��@�U_�XU�UU�N['�(�ԛM�>�pL���0ﶻ�nΧ��g9�^>~+���4�Yzɖ?H��(��1�`�� �S���̫H���qy��H�j���H�(ұ�B�qD�6�d����%��!�v@Iݦ�犒EG��˄z)�6H�6I���@c������(b�$1Ga�&�NV]Ր�B��HsTH���4CT7	�cw���7�Hӌ^4�ǘg�N]�D��-�$�mG�h}.w&@)r��Y�X0�,eA'|���Tl7�9
�Zk�0�c?�s�*�
�J�T�:8� �ĵ^�D�]��B���_���B�.��!��C��8���
�v�Yr��7�jM����~���y�*� q�]�'��-M�����ڻe�GCsF�S>����e�=�6�����W�Y<�ٮ�Ǧvtq�Um�hMPb,T�z2>bw#���#g"G�m���GhF�t�s�/H�kv.�(��g��t�ui�h	&=L�Fl���[�m0��5||*�����c�W�-e��@���C��)�C2��*�0�ʗ�	��[���8ݲ@>����^�c����U���5h�:7�/W�GZ��F;�_��j�K��	�ڋ`wv� �<u�������
�%�<�b�����㪢��d�2��	V�	9���8��qb�;���y|x�c��/lЬKr̹�x��=���i���c�"* E�It�L:b�7���0�8d��������H_����y���g����Z�^k�b���H9��3�E)��lEf��E?���|2),/GNMI��+r��!��$Q�����v�Y4<�Z���A��[�z.�q������cHBT����������Ű9G�HQ��pϏ	�o��P�����F���w���Ü9E6��^p�uӐ��Im�fUK3��e�+�p|���α�d���#;�([�y#3��,0'.A�_�A�#�rp)���zg�T����x<J*�HHHXS�ñ��-�%��D���XVܹ�d�k�FSZRm{)>/SSõ�S�_ڕ�z�rb�9!��j��
4f ����(�Q�4�]�Q
���v{�ǹ����`�prrr��\P�p�Ǘ��U�Vu�pG� �-��~�퓻���84e[U=��D~�*��:��l���x
�2((_�`Ǩ��Y�>8���$h ��j!V���\��?κw�Ha�Z<;g/��μNi%4)�c��}�֞��!�(D1��E���vL�۫�����`�$����ضO����΃EL�v��2%�J�"i=����v*�r��L��vE��b���R�+C�K$�&3�b\��4P��E�Onشn �8�p<�p�v%�c��f�6�U�v��[J��W:��K]O~ą��`�F�k��]���ZH���:�
/EYZ�p��#1�P�f:ȕ.~�M��Y�=.��5��:��Zn�m��5h�W:�]��tݣ2�ȑ�ͳ��Ȕ�Ҕ��M8)[r��v$���&B��H1A�PK�W�a���}cϜ�j�����j<��X�
�� R+�d ���QN,�rѭ�_����)!���YM`�˕��
N���p��~�~�eU��Pg�����������
h�*1�!!���h$� 6�|��{����3^��S��l�̘���t�t9�g�\��?
Y��[r�.]�\#�p�Ԗ�Z�_��G�T^>ݺ_-9/ֳi�rΊ�.b~Jg(�f%�����V�A/"�;���.�o	��	{�OE�;#Y\��}�s�wp >=Y���̑J�z�f50�Ŀsң��Ĥ��.��I�2�`�!��Ot��Ń܂�Z����ĸ�+{�ͯ;�q+m�V��A�����LA�ioZ�o���ϕ/v�Dk�ü_}�U��
�����mA!�e9�Ƌ�eǹ�aQ�Np-�|�2��޽<c�O�+��'Lv��$�]�p�4a���:6FQ��H�L����d��Ý72��b��ӫ�|�b.���4�b���?F�Dɽ�G�̙c�"���V%���է��
�����m��N���+�.��?�/|�Og�͡�MŽ>M�J��P���71T=D�U35Ԓ� �Uĕ�K�:0XM{�pXD�~�)�q�*�_vO���e��|���Tp�h�\�!��v��/D;�>�}L�B�E|��â��{�һU,O{�"����Y_ �!�ڃƌ���k%͎k_jjX���Q)q���0����F0�E/�k^�x�� zT-1mQ��]��C\��'��&�<�e�x��W箼����>���c%}-�~Yw��,�!�����Q��-����C}�BI��B��C%��!P�OR�,������_#�J#<��tb�/X��r�7��Ǡ��͉�A��(�o �	E��O��"����Hhߚ�^����'����D��ч���;�5!�y:E�V�hݨ�~e��bzu�� �Nl$����J��VY�	�u�
W�3͐(���C�?� R�P�����Vx΀@o��Lv?�py�$FE�n������ZUG����DQ�>�ȓs�Ǳ.�2a�|_�jV1�TȢ!'�9�RtJ�gH�;g�Mo������Z �A�G�>�wR��K���E����*����լ��9���@���g͵�����ca��Sܮy��/�~jٟ���x�榚�� �ؤ�Gl��v(\n+
;�$̩	s���5u�{H!�N'�I�z:�d��_Ʊn*��M�u�z�"�y2\fsl�Iԟ�|s'�F�i#���wEzBm��F��S>
:%Q�j�u6)Ɯ*�!��Zܴ�>�f�V���rYL�gw��k�cQ�b6��t�XxtBv��Q����u=��O��Z�|����ш�R)�I�������K�H�`8��Uή �:��`/f<��A�Ge|����D����2���,FU�y6u$�Ͳ������*��Ԇ�� ���>��4#�۹�Z9�(<U�%F�*{`F�K_6�GT�RL7f������Q6Kp0�ZJ)Zq�NV|����e2����ܜ��a�1���y���f�
��PA�P`�X��t;��F��C�W�Jĝo�p�N4�qU�7,�����vb���n�g�����x���"�Qp�qb.I��g/)�ɩP0]п|�0��f�m�)�YZ��v�R!c�M�׿#����X���3P�ۋ�G:Qs�9x^���!�L�M���}�f%��Ǒ��D}u�N���aV�fG��ocV$a����y~jV/�
еl��*j��摯[m�w|���3`=���+����E�`��d�GCÀ&�C<�?��D`8�l���㐒��y/���G�
���ZC2�2�#�lU�5P�4���pi~�25��E��h�QRP�b�}��;(�QfT<�+ ����$lk����EӒK�x���U<�g<&�$�_S�vLat��l�.�9d����c96�1�����Y����*�ga���'/�����|d��#����e�_�QL_J�-�t����N�\�`��|v(AV��h3�(��!�A�'d�O��5�b��N�i��u\�KV�f1ɍ�S���*k�:KAm3�B���Z������G{�����z2�5"&j/oԁ�\/�鰋�*��w!r+��cɒlU;�������s���D�*9��a@�$�(��օ�K~�(ˌ�Q�H�d�7�J����u� L��(���;mh7cLr9���|��%������!�'��׶�=�ٻv�!E�t"ء�v��N�7��gJ'�}.j�;7z��������q@� ��s�s����Rk4
�Lpr�۔���i�aDT����GIǄZ���p�̕��`--��Sq��q�ל.���h7k�VDڐO�jR?��D�����&�kT�~;��ѕ���A���7�r$~�=�'��f�;]<"�[� ��Ux?�d��[�_@�� r�]�ʊ>alW�6�m �����K�L�fe�:�vB(�������y��)�)IFpXbA9.�G��buǔphp0���I.D=ceH��:���zb�6��Hz�?~�yr�H�:�»_��<�6dp�Z��C3���O����#�*�/�Ŋж���~5�t�3_�a�'ś
�x��x��.�fP��o)~���@����Fq9p�����"�{pyf0�+���|�G��!�p���v��V,��o�T��v��/�vkB����:�az��j%Op"�R�R1L�򰰇�U�'��B�)!E@.R�nĄ����)�*}a��e�$,i����'%3��\㩑��}��L1�]�/k<�G?��:1ޕ��}q�^��	Kfk��]�'ၢ��lC"my�sy�q�D�ǒu�H���z���n�|�ü7�Q��r�������p�e+�8�)u�]^��_F�I�`!��bWr^��<���9X����[�n5|E0���_�H��W:�^��\��/�����Ntr?��V&�cN��H���8��Bl�	�(�l7Fa�{��?u��I���/�������r��}O��[�9q6��3��N�D���"TL@�Q1FbJ�C�RC9��Y��Y�UG2�dQ
[m�ӱ��"	¡�7�������*U/����&�D�~�8'1�O�1� F<���\��.�9���`�������^�#�X;9T>:���ů���n�_ڤ�A�MZ�����Fw��gG�S���or>B Z����������D�ϔv�MoY�_��m�R_c�?lr�'�H�t��(p_�l1��Ь�]�_����<����唣i�B\�}�d�1��B��	��&�li�E�����iWd�d�S6��S�u�(�F�ى.n�����ϗNt*X��c���4#Q�8�I�V�Am��J�8[�Qܪ�o�7��d,���V�i�f���0қ�Έ���9K۰ޏ�hG��`L
8��%}�ŭ�"��*�k�5Zh����wlnK���L��2����D�̛�nqq�w��Z�_��ǅ�~��P��8��ݦ|�C���o�������Q w�6��V���Y�_�e��'%�ry�8�K]O?�a
$>����v컳,������i��q�;��X����_�/������g���pR�m%���4�c� "B#�
v����| {�8z��L;�YiFN�H�S�C��4P����%mF�HөF����5Gy�����O���҇��LP��Z8�n�b��P������$�R��ۮN�(�}B��>��]�JÌ�d_B��姚����{��,�3C�'&����ʄR�ѣ�2*���}��s�V8Ҩ��l^��(g�߁��S��jw;�3;N�� ��+�rݐ�-���B��(��2_�T����F斿#�~�d"1�;�/M��PήR�݃ϣ���i����5s��$�ިE>�f��"�f.��44/;����ypE��g5���_%���2���dN���\���4o��2�@���T�YvK�.�8��&��	sv+��q�] ��H��)
�����J�v�u��e	r
�Yt�w�dU��$�0����� �;�}`�9�in܆[$g�����)'����q"vi���>�ׯa��!��x�!j�� ��2F�.Y�T��0I=��A�i]p4p��g�D��2%���x���СZ�cJ�U`{�+'W���/Թ���n((�xj��F�)R��xR�z���vK����Ri,�MqkęounE�L�`�����h��K[��~C$ްHK�U�\8��a�\��f��0�TF��f5�X�F{���D`����(���N(`o���K���v�Z�MQ��|G�u��Y2�(˓�І6-l)j�?Qt?�?�e,嚯�7�X���a�s��� w���Y���wM�����K�$�I~����N�a�Z4�4ɯ%$�
����8��s��D_*2��~B�Ի��&$�I�8�v�`�E#�.��N�P��%UePV��r4oE��s���;�E>�mV��aE�(�j����St�نT~JbK+ĥ3/�OF<mҌ.���0��������E�}�Ӱn�\A��l���!�]�+�,��xN��4�AJ&�4��:�!9s��)�yC�8�'g&�����d��H4�W�E�KC���񯮠7�quue�쌁E�j�gPϟ0fq��HJ��5E��(�_�����D�>�&ueJo�0z�M�.�4y{`o�'��C2�+��=�)x�
'����K<(�r�l�Ԕ:.?�}��7��s9���'D���33�~�.���ϧW���I�7gۘ)	/��	�rG��$(c6�K�E%&��H$�iK*/o]ks��7���8z�o�|W��uq>�?B�2��H�5ޝ��=�Q����]�]O����pzS�<I6��	��fq���rdʺ%窠�.�H��ڎ #����+���s���t��<�VXo�YQJs���%SO,�;
:�ykh�Nر����Z��Y;���ȻU���O��Ω�\��;�t�";��S����V��nN���Vc�T��:�~�A����������T�V�=�	�Bʯ����k��5l�c�E��E~V]Y��)�0�������Z�S�Bgi;mX~�7�ԇ��e�MP�Z�U����.)�&�W�S�����H���bP&�d��>�#���gpw��3��w����kd�;�<E�-���u,Ǻ�א����wy߆�}~f�?p� sW�����S�g��˽U�۵�Mv�<�&}?���$��OsU"?�?�m�Z	6!L���{�o|��܊�ی��fIk�R���iWӳʷ� Oc��)[�bv����x�P��s"2���[�>KdO�X�δ�Y�T �n�<�l8J�&�bT�u$2W9d���i(�	�]����� ���Ɗ,��\3S��y
!ݓ9u�ChUwT���q���^[�ר��;?��P�8�S�z�3����d��^ߝ;{��o��9h��T1T¢T�4v��������`�e��Q)`O /_cа'�v�/g���4k���_�����>{�e����/c���Š�CQ�i����r�ބH-8ܒ����V��&Ft�a1��b>���1�2�'M����?�Ă�&��r���7Ɯ�ٱ�AS�]�g-��_��9PpH��Va~%�Gs�5�0M������ܾ����rSGO�
�(�vO3��� ��3���luAU�f;AW�ϝM�b��.]��ܮѻ�pu�-�6	�w��h�l4���z�r��b�ꐕּ{�-�� �Cشٗ��߷B��@�ݠJr�D.)9;T�������>4�����۟��A1�����ŀ�#���du�߮��jV������!�����{�@�J^d�
���E��־J��.
�+�_��.�^Q�A�!P{����|�����
�[��MCM�ƀp0��5�r��-�v?QeD��sA�rW�L�XAv��6jO0CTq�I*�}
���U�L�����Rt�����d��u����J����4�F�`��7&��,grs�T7��n���} ��C�����,U��H`���X�����O��ѝ0�ާ�+������-mv3�'���8�B�,��e�?/�MUf�ݲ���x�K�Y�P9���e�aA�Z]��X�N���G��D�����o����H��B�� jgZ��Z
C��| ��O Y���;��n�E���zN��3T�N�i�Zp�ł>���C�MI7��w}!����jF�X�~�`���� 'L � R�Y/r]�g�tQ�eS���(~W�my9e;{�o���NPf�AG���l�1j���H�����N��J�̥�Ϙ��M�P+�N�~#I�	M�rᶍ�d�
��!�h�;X�(�9U�h���~u��vk��#5�]�cנ�]6�Ҏrp۾�^���Q�!)���S� RRb�#���ϒ�T�(�U��=����s��Z�c��g���d�q�S��Sb�=�����T��6n�����R�aɠR��_臨�Oa�==y�D.�nnnA.sO�E_�
�#�'��lϑnD�{��j�e�X�?�S{�|X3�:���N�(��>]�<����ɗ��ᷱ��viW�K��Le��� _M̩��{����`�A�P��t5'�ٴ\0FȒ��b��ݿڀ�Rh�_n:3�K?���7�YN���Ӆ�*83����7�Ӯ�hlܚ=x���W&��Z��A��<�-�x�����qB�@�ȅ��	cV�N��MSB_�3�ϩ�I!�2:�W��/s�
���Ň��^�՚_E�0fqFP�3���kd+�k�y�,��aJ�u#m޶�%/:�!y�M�>�u�#����
.:9q��GPaL��?�E���P�f�@��N�����W��חSާ�>��hz���|�	�R8��G�.(_�)��j^+�p��d�;�48H�(#���$W���%���۔J�9/q3�Mmk�� >m���dd��(��,���hJ�U��CQ̹E ��#�M�a�OǱ^��@����-=A@30!b18���3x�.�$3�-pg�%�ی<�Q�S�F�w�e7��m-���
���y��/Jx���4��8�3j�W,�LV-���W�qZ�����gSu���I������-|s�R��P9؝�5��:�(LEyr�h�Eo�G�Æ�B��L�]/`U�����$tN�q�}��tFf'G"�m���u1R**�G/��C����8ʀؖ_(N@� i��5[�:_;@G��"`�PA�%�����-u^��^,*�٠nV#=	I�*���,�d��d�X��1��������H��A��Rq�R!G�y~1�o��Sq��/��%��o4MD`BJ��BY�0[`�I4;�NV�$k~ v���L�|����kt,����14�gPM�����?�9ϔI��n־>m�oo�f��Ͼ����U��Ѭ�Hm� ����J*D����>��d�^�~zR�حև'�{�11D1��)\�ƛ�/�hZ������[_�4����9�/	��č���1�A8ly����F6����D��C� b|�V�P��p
Ƭ�� APq���A�\����d����E�:�XH�IF���
�b�Nh\\�WRI�s��ӕ=X��?����~��)�:4LBD.d�  |N/�>%�A����J����G��D�x���.�AD��P���ۼ�8�yD������E����
d3��y�Z�/��t���bb�����MN*b�{���}K�]��
&n�������'�'���g;4�bK���v���J|j��rT�T�Ӻ(��.2B��)2l�_�b�&ǵ�Xi�=N�6IJ,x�[4�^l"�q��,M��6��#��(8����;�f-�5e?�0`���kVi�s�a�K�8C��������z�!Q���1���Gx �T��:1Q��c��X�0Aۮ�Y�v���>%�g�B��]Q��% ���hKz3�����c�XV����|l�_�FuZɉ�7��k^��oH?lQ��|��|G�0O���U;��x?�8x̝��7��vJ{�Y��>�p�ĸ��)			�m�ߚ_~�SF����^g���k ��U�� ��w���G�/g�����Dˎ<���/ݬ��ILD�(~�4����0����"��d��7����YI&G�c�fS��+o�Ŏx�uzy	p���"֑ 4����@�Q�����ڲBB1,?��_Qhv����p�9�p�����CO��Ή���ߚ�9����'�X�v���n�}y��%HZ^��a	i���y��6>c���������)��1Ѷ�.T?�x�KC�G�M�]��tkb�۶o��}csb۶&�m۶'��v�f��}�:��Z��{�����]]��%������(J0�]�{�A[Í뚁	���W�~:BZ�z��H��/%,&G�Ȩ�r�σ���n�a�=�W�w��$��y��Ը���#��0��Ax�{:X6x��D2�Hd=|���¾���c��a�b�܉��7;,)���p�(�j��Z���0I�����f�}����Q��SS�O�_����l7Z������#�e�Z�cIC[D�rA�yH��lVC5xbIy>eo!��u�8�X9EY0����a�����@�X(��D��i��η�Y9=�4P-����������r��o����2JH�n¬�e7�L*�	ů.J(.�a�-���˶*g!�hϔP�M{�K�vt�[Q���6�[�Uy�Ryr�o�
5=[D�g��?������5럯,��f����
������!}\6lzKm�'�F~�9��Fj�UJ?v�| V�U�w�K�H��ՓY�%b�JP��gh�5��.���J�;W!�����
�+gּ�[[�P��9NQBn����8�q|��U���*���;{7����]y?y��ǟ\���끓W�)N}]���ᓢS�29�T�^p<�F �0�n�(bHR9�:Z������ ��*�ۂ��W&)��M�2n[e�Ev"5�<�մ�d6'��Ѵpw�$2ĵ���:���ɯ~blj3��̽,S(�D�G��x@Q��2��.he���P��<����)�3�N���JQ#R��_���{��� H��&�\�ϮR���P��0'�Q�Z��/Pࢳ��ƬT��MVXݮwOu.gjRV9\��!~�@e�BO:������'$�u.ړ�b��m@�(`�
�I�%I}T�@�P�5�rAI	�2���y�i��� �$ 9I/ο2���##�i.��|-˲f��2IV�!Z�� �bntA�C�FU>v��I�����!�qE�y|o�/	����N7�f���"fʤ	pT�^Xv٦A��2�_!���P	�<T�{��aI~��<ǂЍN�6dS��$xV,rPo�?5�aɯA���{G�rW�����z�z�v�S[_�SB�����z�~�[`�?�kc��i@�˜��-=S�L݌��Y0_�G��Z7�G������"������X���Đ��o"B3+�Øf��o�
�~�Ǹ	>�i��|�������i�f�l��D|\��$���t5X	��~��av'G[�XNס�_v(�Woq"K�z�F0���t����z���(3Oi'ȇj��Sl:�Ku�{�ejC�,�~�\���a�*[����MNb9���m7�����,�6֝cH�B�"�L��5�O{��[#�����Ќ<��%�hh��0?>�Dt���D0_�[1�����l^� O=�v/q1�9�2� S�~i��7���1~���L��a��[�Bf6V�G��Ǚ~AM�������ֆ��
.V_k��O��ɔ5}G��c���s{��������p@b��w�>�PhL���u�A� �C+��/Mj�!`s�m[u��b�:��&� ���6?5���oԓ"4���B��Z�q�l6J�~�8�_8�
t�N7�� u3�q�Z�7��Xc=S����vE��>�%�3_��Yn�̍�vF�_�T0k�+�r=��A�{�ƎU�޲.v#�@�ʹp�W6�VXa�����ص��
�l�f�iE/r۱�4Ġ���9����Nq3�JUj�[���|)3�����Cp�U���7���wX�D넌,��>����T6� N�+�a5ׇ�5�S�ü�D�O7��^��wΚy�Z�^�~�d�j�����Y����W��~�z�,��p�b'P �T��X���
A�"@�)��9J9���Q��{��1RL�jY�'d#o��y�D�4}�.����ڣ{7��#��z8�I(�s�0��9��N(1�0�����A���/>V�o�����f���P9u�H��Y�o�.�(�CL	$/!q=m�����CD�2�MѪUA4�6y��	(%F��Xsǔnr+����eok��9�عKʏ�{���PO��?��_���8�e��۰\��XLG���`�����T�	�//��,7C��g�U���%��t,���uF�I����fƉW���^�2g,G�<!�#U�3��$�R!#qa��0פ\�0�(C�H�����Ć�J�`�	��D���������qd��B����\��^T���=i#,�-�;c`鱫~�X��zڨ.P3�H�){x�r�r�:���Hvę����T15��������\��������G�>��f�v�Y7�S�m�̓�h�FP�e?�e-��I�W
�L�Ց�;>y*��~&�ɝʁ�Y�w�5���`蝓$�8��.�ߞ� 4bZ�.X��q+�#�w��{:l��&5D�$M$Z���xJ�������"�5Y�6/�
��aQ�WC��(�����X�G�o��V��ʖ®��+�RA��3���'��*��FgI��E��?ʋ��͖�$�8���-]��\#��~��F!���@m��q�yuyh{��R� ���Di�	�@�B�W�j���4]L�8�b���|شS5�^�
C�5]�_�n��C$>�=&�A��Z��f�50��!Ґ�e<I��!#r	�����B�	�3�F�BR*rb�*H������M$�۬V߰�7����������Z��X��vf����o|�;8�!�a:�2���A��b|?K|��%�s.xRi���a×��m�ڭoMJ
G!�٣WQkz�%�S������Axx���	�zO�YN�k���_���RT��?���_�[�^����ʮv�*a}}#IQP@�s��v���q9[rI.l��H#5��W�Jt�1�^V��X�b\CR�7��6�Êw��j�����a���	�e���u��f�++��^L���J�i:A����=����/�����)��܀���u��5�}y�h�EC�X���4��Y������	l����=�
֚�U��g��u�,�A��cmI�I-{��F˓��I�t�2.��n2JiAVPA���,Yɺ���̕�����{��oȷgSc����Q���w����P���8LlD/���}�����0|���N�]Lp(�J?�u���yu\�ҳh �ƮW�@Ht���"�	1�׵pX>���e4�����/)�a8Bt��]��
h.�]!!��	|3Ѐ�� �9��K����v�t�9K�Lb?��v��-'5BQ˽[n�6����"��=q�
��(��1�Yk��A9{�\x�֖A�b����O1\$�_kY�\r2������i�	��նMu�����(pp�}��a�ʊ�� ӣ�����x<�=�ޤ��o����+�p�����*��I��HՓ�-c-�'S�^/�7Zi]��$e%�#,��ԁ��_oZ�o %��>���#(�`�Z6x�oI���`��Ci�B���SK�����~�XR�&b\�������;�F�2��������a,�l԰��[b�+Y�\L1���1�����������`�<Ȱ�f���@dW��_��^gN.�Dw����$�6�����VgGz`	$��i>˖.���U�
��Zb��y�U=Q�w.���F9�y��N3�x���#xL�i1���Q�aEQş��p�k���+R��2^D��;�ML@ -����B/��r��&��^�ei��}��(5�r�A&��DQ*�R?����"�9��E�M�n^��C�-���A8�|`i�*�^�1c�	���'{{A��ivgG��yClм	^�!�P�0 �_'?4��PoAfP|�G������8����~;�`@��W�M(J�[��"�� 	��"��v<�����!c/��~���h
�?��a��1�鬶مR���壙��Dn�����j������S�]�Nu!�@�El/It�(��r�1��uXQ�<���}�9�ΓR���~$c;^&��U&δ	��z��N����抱p<+������C��ٶ:G�E���.1R��ph�ꛠ�g�t|v_��<�?����u��\SeNF��4�j��Jr�n'�/���ԋ�6�iW�i]U�ɔ��X�M�q�[l��m6j���gt�q�B	���<�1����v��r��%�x�փ	�)wڊ��4���B CK��%C�@d��y*nG\�%ǝ��DS��_̤#�$B�r�w�T$�۷���n����H�}.��,�n�%���,�L�
�(^���^�-�&?Xc
��y��M�kx�*	��i��./C� Z_�3ΪZ��@�g���&�z������	���
�es��V��&!<G�D�CJUiV[E'��;?N�8��s����j���t�N>�t����%<��d���~r����i�
��y��׉yP{�U͍P�J�u����Qk�_6�?��56'i� Z��B�'N����l�2��[�
�ӱ��P�M|���S���
4(�C�QEb�I�G�!.���,�I1�/�%���V�w�hy)�A���Q��BU����aK���=$�t^�s���"�8^!��Ed��qv�䍝��7}�1�#h��7o�[<0Z
�+�k�?ƶ�l���ǈ�����}�&$�������d��$;��{�Tm�X�dֆ�h��2�%�;�E��P$��[�>�Ы���xxn�Wz@���ڞSk��� ,�'tβ� �9���1R��=D]�~X��*�?<3$r3�����N�@�����Z2����յ��}�A~���r��JK<�u�K��P
��M� ;[�Ň����Wܬq�Evwٹ�ϥS�@��/t�P�i-mq����t}��Lztw(����	cJF��u܌�����h��h�r���z7u��iß��I�iY6-���d��,����?I"4��o��d�?
tvV�<b:(-���W�Y4���V���5s����ݤ�p���D�h�q.!��o�G&�[�����$��;.\V�)
3��^��܏�k�6�R�Vt8��!r��a+��h�vӽ2{Gү�(���A���qC��0�,�p_?]Vrs}���G�5��FW��V+��~>ʋ�	6�~��xJ''Փ_Hy�����~����1�H���x2-����#�n��"�o����<E��.�v�E��D�`6Q<ޥk!�2���ٿ��}�����(8���ߩ��kb�ѷ�K��m\�	�x��� ����)Y3��O#�:������w�>}}�u�h�1��O�)lW2��>-Z��Q��dz�S���d�ͮ��pD��p�����Z�Ӝ`RIBA,Yb0�x��|�TQ�����amu|=/����3,��攇M⵪�H��k�*�Z:��9�E�q��_��rQ_2+&��X��s��=���̣(9ÆWb��-3u$@xƜ�$ěҪt�BzHPɨ�;��gX�U�G]�fç2�w3�����K,�^�#5,�(���	�`g����m4�����k���꾱��%��)3E��:��ris8ۀx<���r���iKfo���	ϸ�{�a�K��L[(�#a2�8���ٲ�*!�x;4D��G� �������I� !�
\y���T*��������6Ȟ�??9�X�|��Sړ��,[Ճ��)��Ą�d8�%UY^t�B%�P��-5��vG�⓶L���>/����
���"��nqK�q��u�<Ko���R�"�]	�b$��XEa����Q9�]9Nwl��{axP�뼋��seSVk��\�+Q�˔] �(K�s��a[2��?�w�-Eж����o�d��1f<���r󦀊o�V6�?�X&R���;�PR"O�.D�DB�[�)�ؘ�bY���������8�~�"��U�Z��`���U����t�t�e�ߑY��(�OY+�V�Ît�0"l�$��i�b�ns8��O�CX�R��f��J͆�7YS���?��-����"bJ�/5�G�>��q3�L�t�=��;�'!� �c��/?��5��6�2.��)"����7����
pih�Z�H�  40�{'��;�`��߸I�'[M?DEɃ���L�!<<~��0��C�>���������O��e)GHY�uYQ�|��<}�T5(�ga��.~E�\�����m.'�$���fN7��)���h�l����X��G��t9��y��c^fD����4���@�׼cT��`�R��������v�q��b�PXZQ��u����5k{��d����T�|��.�k�>�F�P�����7ʈ������?R�тU�G��u;�z�~v}#��f�ż΁��G�O���u�P�쟾o><7?��R�2���<��j�0s�`�ي���訍��v��م���j�D�=����f%�٧LGYx�4��+#���R�����&�:�q<�=/B��8Ȋ�T������� ��%���C+���I�A(\�َYMR-��{Rɕ+�&�zDy��A$��X�ie.�3��v_��cЪ�J
���̳��*/��+O�3���<}����y{~]鎉��%i�j��m�1�-]���K=KU&EE!U�"�[o�e��;�<��'��W"�{��c�2v����)��"�\�������J�̖+5�9cබ��q� �;F�?4-?�+��so5P���r1?h��Aa�X�����^�����~�}Z�ɊYH��8��SB��%�abc3���%��;6�m�D��4�9�E6_U�z�w]��@�@|�$�ʆL�R�؇#pî�������F��{k����oW��ց� �W��,���b���J�p�a�Ӵ;�l���$�rj��T����P���;�A�'ѻ���z��(t
�Z`Bq���|F\ s`���y����Ʈw�27j�፮>J(�V�����x��ds4�O�@�I�t��!����ᛜ��
(�nZu=u����O�!S�W_0<�
s�fx� '����J�n�-)D �26>~%���B����ޚyqr�3�)D6m��{�
�){��y^hq�6a��`l����=XtF�3�����:�z���]� /�2sDH~D�h6#!E�s���@Ԥ��:�U, U߿�'m?r>XL܎���e�`!��=s>��u�i��r<�u�{�H�gW �[�լ��U5H��M��0�''���!H�ׁϻo� ����Y�L,�d�b����q��m'>s�u�
Z:"�A�"<����?� =V8��I.�ߗ�}1!�D��qR�\f �;XysCN���]��#r(�Ð�l��EJ7}�d6A�K�F�F=��}D�e�0��:l�99�*|�� %��g��ӣv��U������ݭ�������G�Pv�7�X#�0"��I'��6'Y�c�\C���y���}�4��!�I�j�͆|������j���-��u�W��!*��$E=t:9?#���$���>n�M�t?}��z�<�,w���B0�:�
Q��)O�H�,?�Ɣ�����h�/�����%E�ְ���I�����@�s�Q�>e�<����W���k���t:+ٔ���]����e��E�U�V,@�P�(L_@hN���p��a��zE~�D�l�ܛ0]��4:�4��h��͜��O�NC&�(�����Z�fϻх������ݮ�`^n��5��ڵ�>�jEK�&a�!�^�Y�k�c��(\-Nn4x���ha�h�.$�L{6.V{�;������z��km(K���$!�c-Wu�D�1��%��81���i�nOT˅�&#��!&��4k��4"u��AV�Nji^���	N��u.�`!��[y�0�8=,�<q:�Md���jD���t�^t������~4��w�}��bF�mh�����g�����
�����G����M{?���ܼbH'�]pO�/�\�EU,�k���({�h�W/�<"��y7L�?�J�y��g�����~�p��"3_`�PܴA2N��E9W�G=Y��G�X?�l����9�N�Z������(ve�����# ��q���YV{�V�p��_#�A �Ve�r����׬\{YE�\�jV!
ŊT �������(�_�b����$�>�*�Ṛ�YTYw��-���W�Θ�$ut��
�s��賣�`/ԧ�5Q���*Uw�w.��MrTF���2IR�� �p��y��j��S���M�F�����Z4�W�DA<�ɺ9��h~�w�*d�3�9f�A�`a���*��k0��6	�E��Fu^S�	rN��́���gՇ��o��6$�#�1�4R�s~��M`�*5��aϝ��>���扨r86M�����>�g��z�?7_�����fƼ/��`I��(��.���/���K+z���9^��j�5N��<O�|t&�Խ �1���{��f4���q'|ç-W"44���YNf��,�5]ԋ�&Z������u&�}�Z$J\��d����9��M8LC�Pz���uI�;we�ϯǂ3�v�?�ȗ�REb���'x6�mOL��,E8^r��X���p|>8}{^�C_�>����mn|o�nߎx>C�M��E�7W �cd��n�˞
b]֗n���&�6���Ix$r�}������%��s���z ��[�A�q�^���!���5�Ϧ�ia�yjՋ�_�
i��#�9�m�Riz��x	/:�7�	�H�yݘ�ۖ�X�ُ��wK��֒Φ�x�6.�+�$���j>ʾ��2[��e�YB^x��X�~+�{lMk6n���Z.ႃ�S鬙l����G�����#2`�P�X����J��<=��~������ʲ�l{���?�C�,u����)���dwB|�Q� �]�:2��]����e��{�~�S�m]=�L͂7	z}����۶�F�)m���l3圁�Y송�8W����[���7Պ_�/֓����Pb1�����*>@�7���Ue������.T�t�!�o�1A�r��{(�;��2������ѽQ<����27>��WN�1��Ua���u�;��]7�:��h�]o6#�x�5qrb^	CV�j�WV�:o����=6�����\]�MZѺ����Ӌ�(,�\t�����������>]�?o{>�� �T��Xg�9�-JƇ��7���U`�ҡ������� mΠ	z&�y`R<^�]mwA�..�C������?Ю��|�$Gq@ᄶ�?�u-�Q�4�L���'���4�^�Y�k��݄S����������o��͜��M�V��}Pr��x!�L��`��5>���ar�Ӷ��q��dD���Ⱦ=�
V����$� ����D��&҆�ǅz�m|j��z:�$k�v_�Pۍ���aS�f����O���.�Qm��C;=�ÄA��.F7ݾf��F�Jە?t��=r��ek�\��Z����5����a�|��evF���cg�~� ���*0�X.*&��h�<m��e�������8r��C����h��ɥ����z�[n�#&�`�2G$ҘC]p��O�N��OqX��p�W����ڀ�H9���VtL�]��5�7rn��T��vc<U8��B���g4�5}��u��o�KA������@��J/���A�``��
56���@�MD�p��	I�YM32Ms���6YMa�8�3,M���9H9*�M�H�℘�H=i=�-=��$x6���F6B��n�[r�8k~���x�g���*�e�hX+ё�
E�s� G��N����b2`j!?�~�P��U���_��� ?�D�[��0wS�5�&Z n2޼�<�{�~T�9G!���0��+!*��
"���>
yR'�ƨ��M���[j0#�����{e�-��C��hr`���J�ZQpq̐?K ـ�-�S6�8$��r������?h�#?��W[�I��G��,�J�Vt��J2K��-�:⚘hJ���z�q���#�)�:��)�b�7�[��e��g����+�F��kZ�X�����;n��H��ً#,&��~�x�����SCDЗ����(:}V��O��O ����G�o%pV'�-�:7�hSx:�L�]߅��6�����f��
�6n5�p&Ҥ�ۦ2vdԞ�C΍�>6U�!+�4%!w<�V�3�a�D����G��sj[P\���&K�a�n�kғh�ʈ�s	p���Z8b��E�+����/�V��Y~Z��6!�^$Cݝ2����s9:+�
�Omx��� n
9��'I����X�@%f��Z���GIn\���e�:J�	�1i,̆���1q��Hoxi���J�0����ΓU����D�CN�
f1?�؁"�g�6y��ْx��C���m��X����9���yڽƏ�ǁ^��ל��8cw��sQ lr�>��5���tc\����X�`�� {��t�&*�k����5RO"�d�^�̿������אC�Ģ��xÓ��[�?��Ͽ���������s�H��Ә�3�v�-Z�t�����_n==C&f��g��s��F�ա�{dc��S�5�o�f4k�-3���ǋ{�^����P��>���.��6���1�Foj�&˅�2h~�� ������h'].
\'�i8�3|���=�����.[��pi�$���>�������-z�l_}��<����-'�v��[e���A�տ@�:�LI����Hm
$�v��l��r�D��=N���
kqM5ZS^��V�0�{,Y��ξU�Yk��EQێt@h�x�2�\L���q�!Q�s�u@0�q��p��֬XR��M����.Տ"���V��~�LD�b���ӹ[`��H������t��Bz�d��S;���YM�?�,i�g�J:�����ɂ�u/�ӭ�6�*B[s�������6��Z�}8�m�a[M�����a���) K��Q��;�v�3�ϖ�t���E�����o�Wĉ���u�&��\߳��b�j��2:�>�Sd�^�$j��|F����2�m�:�*��2�έ~q�x�r�߰�pP��!��^�;���Z�2�U0/�W(�3GGP�a�BItq����)1_O����Ğ�o*�1��Cc�̂��f�~Q���\��i����v�n��W�?;I¼jA'j��0��q�6�[�[@���$�S�4GV��T�*i(�n5ذ!�m�Wi�R�Z]<=D&�=F��Vm���I�C'fx3��ζ\ Ju��Tdo�X��0�F��Ր��eky P6�{߂�Qr��e���C^�x��F9V�x���an�"��7v�}��h��L)�q�n�j���ݵ���K��k8��-�F.�*������2P/�|Ʉ�L1}mrO��Y���ݸn-(��/WWZ�?���aD�3��b�a��f�~�R3kD�aq��7��<�Y!U?ųEl�p{,�#)����;�CV�G��9u*fCM��jk�aG���yǃ���D7���;8�[-ƫ���r-�z��D�����oφ���]��5�[�l�/�Gq芖�sݧ��3*�h�Q܈h�2j��]<cd�O�5��($�ʾ��Q�|Yg�v�(J��a��|���  �!�E8��8�S<r���?՜؄?��W���t>���H)�w��c�'���5?�7�1:>3Ɛ�GZp�1N���r���_Gw@{�`��9>|�� �h����XD7��r6�ѕ��)��KT@��.�CֵpE1�_��;~�S��:xl���j��3�A��{Qۜ�vO��;����=H�g�K��j�Q�xp�G��?_]~���b2�?����!�4�ӎ ۲�šȎ��G�1h�V����2��h�~NU�� =�B��^�o�T����q��q��i�kt��'��+�>�BA�?���
l��Mt@��4���~�;TH���|�*�d 9%~��|f�!�=j`-�!�³Mg�7n�����f��C��.�-��I�Y|=�a���]<��Z�	�^���7@58��?�e٤�mv,R}y��|g�1.Ns�E�}e< h]��xch�.c3M%�;1���ޥ₭��oy��	+Uy.����G���)�8�P�I.]�2��S����!�(�h�H���÷�=��~cYz�0���[_m��e�s� �z�QP���k�Q.T����Mf>FJW`� GfHY��T�̊����,��B�(�'��A����%�ّX�����IU�̙���B�=��uZɡ�0ؖ^���`��?T�i�����EH��S���tE"�(hЈ���0�0iGp��㰖mR�h1��Mj�Ԫ�����?�sd+:����d�;����\�"�̰��S�뽪)"���U]~�����!� ��z��5j�Dn�m�G����Z����z�WfF���猭�&"��<��5�:��H���v8:��qݻg����?M^���=S�e��0s1 �[WI�/c
J# `�39��)�?i-��}ZtK�����������#�@�''�R�L��|�Y�ۮ���[ ������κ� �0���ޙ�bDa�C�ӠQ��i!e�`�X�VT.�4d9B��'�'��h�j�/��ﷶ�v���+��E$4�gc0�I��
��:
�VR�7�5��%>�[vZ3I����]<{�b��������t?ή�icAp�r]�d�\�1��� �܅�%%Xp��ϔ����Œ���������cdi��4��v�ӓ�a�M���yՕ�1�;�a��۷ϰ@��N��Z�m��{W����N�'ONOW�e�^�I�->5l��G�S"���-M���G�׹� u��;pl%�ۺv��?֨fE��S\��O.��c�$U7Ųt0c̃M�,�iH�01JۺU$S��{҆�r&g���SֱY��u�е�36ʩ�x�[�HM�-F����P�X���FB��������� �qH]�a59ӗ@�A~�\o�=�'�SKS��E�p���[�'�ЋB�.s�������Z<���[v@���L��������Wm��r��U�0$s��`�vC	{����շ��O��^5G�M|em�v�Q��~�!C�G���[H^w��T6������">���o����l)JL5�D������k��O���+��i��Ǌ>{o��@7'�8_��E%�$JD�V�g���A��?�������,ޤF^�٫�Mv&q	�󨎯U-DKvrNA#{�YO7����c˴�k|?μ^*���y�����mo)8�KS�r���j�`���zpeyo��O�5e4P�D�Q��I��4�ƶ�5aV�idMM��Pq�=�&$�ߍ���7Y�v�;.5�&�E�w��v�� ��S�����B� `�._t�F|Q=k�i��aT;��"�ϕ.1���Y�-��
���K�_�'^�o<L��|���^�>k�6���EDWS�##ݰ�iu�ɓ�p�];��#�Nh�A�F;V�°�Q(�)��U�{qp@��P���؄+5�#
Ht�����p����-'�Ez�	cR��c�, H"�p4�����;2W����p����&�G	�k�?�{(�B��O�}��e'p\G����B�aE&R���S<���c��'�35Mj�4�;ȝ	Ayl�R�i��fj���1����Qʦ�V��]�	��{{��T�j�~�n7s�T"t�����boq�N�?���b^�Ѥ�JS`�l�FO@�ov��#��KBH8���Id@����a��|$�W�b[#RXs�U(!Xr��&�M,��� +L��5C� �3�
�m�%�R�����j�My���ߕ��@S�]�d���0�b��n�f��f�H?�L���D���/�j�m&w{�X�6q=2��9��v�X��	Ǖ"))�jZW�"���F�� �q�Q-J��P~����Ȱ����A���`j�����Lfe+���9qVhV���8/��]�0���Ms����آ��X�_�%P�,�y�Z���VU�#h�� ��V��N���-���T`���˕r�边��P�*IP$=aK�++'���6*M�;��� E͢�S�CE���+�N��VH��zϠmP_�	��1���q�ÕQ���6r��fם0X��>�d���J����*6ɋ5�ea\���zN&�nI,���BY�UA/�BxM+d��t�$�-�2�|U��^�chZ2�j��7���l�Ε� _��ˆ)6�6��o:�y�ܾM��t��¨���v�e�3�F�+A�G����ٟ����zC��]�P�	EN�rI��#Y�u�Z�i�\p���4Y���?�M�8�׏�flR8��R�^�[���O��� 𠐛���gd�ǊD7L�;g�%��m�=af<�6-�k��N����]��W��#IV"��b���c�uc�	K�e$.CR*�"p{͸���+����h�E�A�p�pE?��D���G"�}J��|�-����y�V�u��/���.*<��\pfb|!��?i���/l.D�j��9{oǍ�l��:�Cf� ���h!�C�jhu���,f~;j��D�z�I,�q�
����(|$�x�@�M�ۇ3���s��b?F�ʤJh�T��FC]
ER ���#Qb�_ x������E�v@����/N���n�~��~lb,H�Ć�� ���>��"�F[6)����t�cXow��+�[��YTe���|=k{9�L�n�M>㼧O��0�G�Ò�K�U*iK��w��ss�>�D��DR0���v��!Y�Z%H" _6+�UnW�GY��-�^�(�����w�w=����U޳����Y��]�Y[��Q1Ü��_�
�k��MF���M����
�����#+5�������ƌ�\�Q'���-�p�\��V�6}6l�^GɼR��޴w��yc�9O���-��2�~��A�%��z����g�6�tm-eGf���(���q���z_p����3$�Ϲn2��{ fǩ����ݚ��� �G�-S!]ʗp۵�W:C*��ZN�>Nbc� �P
^"{��r?ޏ����܍�ܫ�����3�D4�i�R�Q�n:�j��e���I ����Eo]�x&\J�6~�>]n������RS�8r���.��,kp-�6�|�í��҈_�y�9l�߄�����@��+����00A����h����'���*W�(9F�H߯p����o���\�5YI<Ⱦ��z��!����������$���o6��z�Va�(�Һ*�X��3��Ei�0Ɏ�.T?lD݄�*L����q�䶱��B���P��O�h�����S����A�
u�7w]R�l���<���Y����T��P�%J?h>�B;L�nT���>��?�؎9ĢYI�������;N�#T�e�D��[�����|��R�%��@�ΡJuAw��V�U�!uR�5��vl AЦ�A�SXv�S{�$.s���!�S���<k;�n��� x.�;aФuHRN��+B���H��j�k��Mn�����*�v����IAS����<�j�\E7S\4��t\�o�����B����ې}j�/X�ҙOD�/?���kcdۏ(�'��udE��w��~�����E���.��M;�u`�Y��{�i��L�G"���a�9#��M�"�s���_��G�Ӏc�b�HJ���������B�`j!����������R
�(�z�*�A���*�Ũ��"I
"%���0��s�G�g�B$����@K�!��H��9	��h�Ȧ��נ�i:��&���᳟�G�$;��IN�lK�'��?��z�Y�J���S��4e_lKSf�; �.�� �Qw'��$�HG�g��Q�5K
c��a�)��~��)sF�W�&��2�fe�Wy���|��b}��>���)j*{5���XTW?�?m��u��Q?o�5��zc�;G��!�	�F�������l���<��J!�a��aB$�����5��E�Yʺ��cإGJ��Կ5ots�* �,(��£HcL9i��YU��q��fߞ��SǴ��7���1�tBY7�b�C���_�-�\��m�2�p0�"2��^��p$@'wΝ��H�!{tql��H����P�ne���?�������5�
u:���zQ'��D�<0����S39^	su��ݯ��w�3�yR)��TsL��G���IHJ`�$�˘�MB��F����I���)S��R���A�ﲯ��D�"�X2G��k��6U��6�[}��?��1��.�F�/�8y�m۶m��ض���tlv:�c��$߬���u�=�]{שS5<��waN��]A�X:�t�7�u��CPXNɽ�3�k��n�~stt�2T	��Xr����Ɩ�X����sƹ䠱�J�1u*K޵͔�� wh� ��8�V���q?��6E�nk�j�4�n�Z�)F,8�`�炎�Y�=kZ+%�Af���b���r�vC�Zm��Dx���{t|y��i�·ߕ�jl[����%��5���z���%���b6�9R$|�_2��z-r��R��|X���U�?���կ�'��y��G�ʔ|`(g�[��q�p�X��)ފT�8	�0k�`h�ޜ��w��Q�$T)��Jm�+���rX�Jf�N����o��Eۙ{7٭w`�%ů�u���2�9z���c.v�|>�����N��}�־O�� 2�����b�}}3�+����N�K
��|�^Aq9oW��Y��ʃ/U
l�P���3%��{�N�r�*c�߀װ�xDPohl�ܫ�O���)TQ�4�����4��o����d��#@|P�fk�Vu=&�ѻ�?�PY�-��`�H�W�y�����)|�'�/�Չ�4.PY/V��OM'��M��1�q/�خ� |<�GTSR*m�� �KFa{�Gn�Ԫ�չ�P`Y�I�3˂�9|&5�@rꇡ��Pן
K�.?����w P?L����������a���:,��08|�k�Ewx�#7mM�l��aq|�ŝ�L��7��I���d(k��쟟�_]�@Ī�T�V�F[l��E鍆"SN�~!EKG� ��&j�̈���O8{�<��c{ws%�C!1�:��{]��ܷv�4��+T�Ŕ�	�]��<�N�����&Z	ha�<e+�#�����L���AJޟ�3gO�ߑB�+<�NZ�T�(�@����'���#`����i4���a?��T1�1�N�zsV��D��Z�;a���`P��.�;9�=�������'Nu�*�.b���n�뾓ڃ�!����ݤ���&Y�F���ٜc�J!�yω�y�����E��	<L�s��_�[�It��h������w\�-v{��\T� ���T(��o$|o�ʔ��+##vk�<� ���5�?n&&ؼ�Qٝ0����dI��)R%O�:������A��Aȋa����g�f] �����62�.+��Ha�H8�-Q���G/`��#6�:��#x��Ldb?�V�Ds�JN|�5`+�,!ǖ�Ⱆ�z3Z���d�0��j�Rg�,,L�����yJڍ�5>��<a�w[����EJ�� K�J����s��^g>C�R|Ń����ll�1���&}b�O�VaG)�9Q{wj)I]��Ǉǹa�Ֆ6դ�⭾Xx��!qp��"����L�vg�ޓ�b�+���H+o�+ۍ}��4^�9%�� �IUH�]�6�Z���K����N�E����P��ޘ��QzztdY� `=�x���q�F���iI�,
�vU��]��D�9�*�vԙ�݆� N5��S vn]m�ҝ�A�۟���\l�r��*�K_�\qd�6��*	
�G`��q�V�� 0L�#i��v��"X�\5� 6~!i�,�t�i�� :��A�x�p4��g��u|��y}	�lC�D��E�d{<��?�$�v?3YWr��E;ԍ��W���T�`��٢�9n_�A`�>$k�c��:�/3�������ݮ���^�O�%"l�$ÄS��賊!�͢����o3El��k̹��fvNbx{����B�n�C�ͻ:����"Q�R�u�_����8�Q�vɷ7�8ܕ>���#Y�E�`�C4�W�us�����R;������c��$��C�7QH1Y��<���	��
cƩD:����s���ǽ8��曎�g����#?�걫x��b�crv��0�c��8ʜ�K����e#�w��i�̶�V�^�e_��ʸ0�Ǔ���'��8,�4��P! ��,�9����͘O�)l��� B�F�T4����L١����&0�rGZ�{�R���]�(��\�D����HZ'�����Q{P��O�r�&�!�1��_�N�J[o=���Ix�VóL��Ї.�̙3�t���]x�*���IT���A��y�"�ʥ9.!�L\��{?fs;o��U#��@#P"���[E��ܶ�����-Bc��}��(���Y���,R
n�:�:��
�Ly�;tCH&�3�[^�P�UT��E+�O|��т���-��8m�B������{y=X��Zo�.�p��"��a�Y�p��;��(��
��n
�ӓs�P���'<))�{����9ww�1��Q�y�7"�7���x�\���

�	����1[!kZEN���Pi�s�)r-CCd�څ���V����GSz���܂ qEdH�������&w��pJ��4X�5���P�rYis��}L�ʼܑ��<�����r��L���{��]uξ��"v�����ƮV��OM�ߘ%�nڎJ��.6�+Ti��j
�?�ϥ�ڷ:x��`I�39L��e���d��W".��>INRi�k�vS{�C|��k�-����������Y}]�/N�dp� �HH�Td��J˒�ub��aj��4��q~�6����d�:��m?ez?Ŀ��V��*=&�x_�'�݉I�W��'�g�R�.��Ƒ�WYTb�Ӄq&����g����P��5���'�-y�9N��� ��Xj��N`��o�P�:�6�M)=YM�}�� �2r9K�U��<ϕ��k��X��Г�}�k��Nm|���Z�R=��G!�2d���9��0]g�F�irZ*s��:/�Azգvլ�=���ѳ������-�v�U���6�2����>dS�!%�)n�TcZ�Hd�i�H�MKr�Eu:i�~�&F4�t���l��4���ח��qY��7g��)���ʧ�Y	sD���soㅆe�ɧiŷ-~�U	�"tt62P��]��j����́�ŷ,�"c�[V�{*�Lz�w�&��H�����U�vp��M�|��,F	������-@�J�"��! 9�$�v�UgF]:۸Q��ѱ@f�����W)G���J��5�T�7Q=Qrpꙓ���Ś{�"��=`6je0-ŕ�.f�0Fn@"rt�f��B� R8M���~2�5�`�?)����ѿ<.��/z^�	J5hڞ�K�z��E��1֋���x��6���v������؂���������^#3L��m#E�J�8���D�l��Xw�&<�aX� Ы519	o�n�/����33=ǔ�Dz����|�@�` ����R�{aJ�T�v��ǣ˛�wr�҅�ig,ϝG�� yRXLM\����mx����k�ȯL�{��Em�3�Yʑ�3c
�KЅ�p�s:{+7��xeO���Z����o�����e�W��_�J>6��:�_�?,y\w�C]���4�Ѣ����%B��a\�H�Lﴯ��MM��p���%D����`�5в~�%��B�W���P9�jD"��� �w��&���$.Z�Gӹ舰���T0����]ۖP�C��UL-:5Fav�� ߴ��:#kP�]i;?"�d�� OWV2#����$�.`���T�-=]����0�Of_g��v��g��ϾRm���qQǉC�P�Y�s;o%��D�B�#����oo�w�;y��r�`س4�{y�$T���-��2̽�$�q��i)צ��kB""9������qW�'�ڗ%v��>D���Y�1*@ &pa�ճs��'6�4��ݱ�u���I���6��>���G���Дk�hK&��Q��.e܀N��2��|���$!���U�����v��=��p�_����O���,	�	��y�Y�u��ɋt;sG&���3!�x�`��H�}j}ά5� '�dڬ�?1W��I~�m���ֵ9�F�ٞ5�����g��"�9O�[�Z>A|�����)T=rG�[��k>���"����e���9g<?���y��~��EM��dW��0�L,��ao����4��Q;��g]k���Fk
ʸ%=?΋�]w��I��{�'$����B�m`�Q����7 Y#z����P"�%�$}C6L7E@IJ؞�^8��d�qU%2�x�=�e<"�|�F��2aL��ḻ��	Ct�B%�����A������JY%-nx�)=��"̣V������A�|��������9�u�g�m��y�ٍK��H��g?�|4�m��o�)�{ޮ�!A��h�0��VF�7037�
��#���n7|
VՍ�X�I��}
h0
���W�����N"l�8�X2�Î�Y�gI�u���A�j�z�?�8O��c�\��n}�7��_ېn���=j��,���� �r����!����`gglA/�W���@9LW���1}	f��9��C�5)����SŚ� Ux�sW�z�F�^ �02>�z��լ��c�v��ems�r���qThp�F`�Mdmh��U����W���Rv�0�~�A�GB]"��GU�c.^�� ������Q*������iv�1 �B�MG7������EQ_�K	���J]f"l���Z��i{��Z��:���>f�Ҟ��׍�q��.)C�w���[b��[Čۑ��`K�˽�����f�ܦ����@���ٽ��sw�=��k�����ޛ
|���+cyHK�~��:�Wڊ���@J+4�'^��Qֽ0ķ��i��[��8K��t�pmŔ2�l�l۬���n6��O+�j�[����YzA��V7�8�A7S.xx�ȬQT"k���Xf3f���7�.5�AJ��A�R{ȁg�#�4���®�`��!z�G�� �4ߋ�Y|�渴js*C��{� IOP4(CJ"�����ϻ�lV�K2�Kr�V"U6�[�r5�-I.�T#7��y����*X^|��2���lG0��L�SgL�0��hq�A(�F�FڤINt�81���M�h꺮�yΈ|[�Hh�����N3��۵����׵?��M�tA3&	��dS��ж�9M2�(1��O��9	,ZzBƑ�Z�Fy�x�%J��2���kg7�qa�Q�3�5'3�{��}��uM�T�c2���z��@�+�D�St��l�qZ����AH�~�F#68;��E�j�Ҏ� yaN'Q:����C�T�� .ƾ���Hms���VZ!���8͛�<�%�io��!Tg} w��B�8�@2���Acұ˓�]�����e�(�V��0%3>�fL=�y 4��Q������&O}W<�����"��zuƙ;E��Z����1BQ���t�l!A��"1~A�f����(f�M�h���i΃��g[������%T|\���_����ɲYl��nɈWهd)..���gT�.�L
��t����f�c��D�b'ƾ+Q�D�]�IU�����$�����H��Q��6�|���0_g�y���_1d�=xJ\�+�%a?�5�??Y�݁��^��m��%��e���9�?0��t\�D��i4'r�7�b񹵞�w�on��甦�;zv����:�O�%ipu=����l�T����r������n+�߬���Jl��'s�����u�$���Z�;���O8a/<�;����yA'��\�9��O��wC�Iö��V�[2�!�Y�
� �T,Q]�ڸ�*mk5ǞY�uɔ��NM{���S���^��lm�pY���[3-�1�-	�sN���'�.J��/3���c�I2�s��-�"������˽y�8uK
\�W�!M�;�'3�<�O|�;����K�%4u�iQ�-�"S����Z��㌲����^ݧ��3�H^��/���5��=���L^��Km�2&����꣨��*T!�\/g�T�a�Җ�L("���Ȫ�Vx��ʽ)�^W	�: ��OJ�
����`^$�\T�"��
�l,|�(g!:n	���S�jNYIFMc��,©�m���q??��W,�6����L���8_e�)n�Y\Ywt�BnԔ�<�]�ü�Г@\��Y��h��nw$��ڏB���i����N�y��ܪHGX4����P�զ���~�iL��	��z73�:���T�8ā(H�8r?�[�X*]7��t��� �~Q�1k�6�R�a�-
��t�\@jM+/��
���y�M*i����� \�M�,��f���-q
�[ �ǁ���.�QZҒK<�G�d�G��<�U�N��"��f���j!�#�YMNN^v�}@eɿq�h)��<ブ��</V�5`��k��v:Mq4k���]C��a�9�3�o{����t�Ͼ�5�]���_�Tgdf��w�Ȗټk��'Z?EN�t�_ϑ�bM�E��3�q���mbmh�:n�-�$�i��אm�z.1mx��٣���i�w��;���߃,Ld�s�i�t ӠѢ�Lv�pCH=vU[��0:&��45J�Q���U����8��t������[�r(�_����"�H��
?լZ'�PI�`u�0�hh���}���.Ϭ��|�l��/����'tiM�"Qh��iO�<�(~��"�I�l��̎����̠#.a��pPn5F��Vwt07��0�ضO\]FZ�Q��Q���j�o��v��8 ��g��&���rana�#�y�6���*��1�_@�OL��������&Q��K��YԹ_�-Vi�o�99>��("�y�_�=glQ\��1�
��>^g�9=1*��R���_�ک�� �I3�q�	��A�oa6�w*��;��kA����Q�֋2���E�|O&���ί��fx0�mÓ�P�ƴ����qӘ��T���>��0�am5b�Yf����a	aa.a�2�P���V%:�N*�"G��\y̎i0Cdl�=�0*��(�:42>��w�N��ۮc�Z��v�G�.���~U�AC�T�u'���h� p~�ٹc���i�c��Q���P�x�a�9kz
r�w|� �u�'�t�߱�������0���9zsy���j�2rs�<\�~a���!���+HU(�0����4�b��ʩ�nqX=໸�}��	J,�i^��غf�.�⿊�/�R�^�ov�$G���p���nb���������߇!g��
��q;����8��'&���k��� [_�#(%�m�D]�T×�nMk=������4��:�s����-W�hQeT�w���1��3�~x�:o$.K89�Mr�8�y��PG����|���@t��v��7<��Rd�b�`{Խ��������:�)��F�ɚM*��b��௻�}/�5oIY\���&��p��?�
 c�o�	06�!��p\A���W����w���rO��[��_0i�BL�Ľ�ڔa�Q����hr�5=�C��g\���Ρ:�C>;hy���i��֔(V�u��☏l�ށ��'�~~0���l��,Ml��}��]_
W�Q0vV(M��G\��+!����w7�`3x$=�'��?��R�����<>��{?U��OU��GR(,��hA��������# UT7k��XF�V1��t{�B�k� çK�����C�yγ7z�?�0(V�$F)p|�X;�ɢ�{/_:�&K�-jf��@����d�[-e�5�X�_ɪ��Uo��,P�iu15���h�+c΀%�����w��*P�(6�C��{2F��g���%PF�2�y����Cpܾ$Y��&y���D.��6��u��F���y�t�I��ݎ��#O��N���/	:˥��%�cR�z�|Z��[�P�  ����󻬉��ɍ}P��f�fq�kHb���^^�n�԰\9ݿKvBސ�3P�0����*3�%VDW�g��bcdd�;^�z���,�%Ay�FP��w"�%
ǎ�0�%O��yrU�fQ�KJjG�`lu4$BP�5L�����̯{AW4s|�Ի����~��	�I���y*
�sf��{�y�=X ��;o�Ur�7�'�)S����D%�n�g�����l�8d�iE�_���N%;���TR���"Tϟ�D��-����.g��}�0�wG��P��ֵw��p5�Sn$�&d�_�D��9��ı�śTwT94OÄ�p���IϷ9N3S�L�+�>���儓�ؔ�h\kQ���T��ޛd8{/:<-�B=����iХ�HF�0��^���f�yM��e�i���KRU�vH�O����E��C$H�C1B5Rb� ���^^yrR�x��ff?r�+����A�1���)%R�7�}sr��+F,8�Op�T��Z`N�\�!Y\��3尭� ^GaH�/���jsv������nN��v�N��e�- v�p����~Y��^Ĉ�۠��ߚ��t\����m��ۭ��k���-��F��n����� o��N�5���S�E`��O�D]w�R�9�zH��PU$�F_��1�G�����I�,��P�s��j��  ����Jc@��נҢ�t����'g�'���O�b₟Dod���Waҥ��W�9�E���v%��z��U�\i�e�"�	�_��D�E֫��U��g�� ā+������Xލp�
��qʭ��ce�% [���xr��� Ak�OF`�$���k��"hFM��_��s[��r&�6��]�X[���>;��?���=�O�F�{n�����0��,�S$�\,H����bg5B*s����Jzy�����]�Z�#%Q���z�bD�(�\1���"�Մ��@t�EA�d533�X:����.T�9S�zLXdy6������5p��R���Y�Aq�hN��G8�;Fk=�9a]�֟i1��Ũ}U�u}n�Xl�q��ꏆ"	%��s��
���q^o�뻤��VT��e;?9�xy0��^;Ҫ#��Ʀ4�;N��d�~-Z�������L�>lL�G�P�FiE�q�.�z����>� �ܡq�w�}��G���eCCX���9$J�)��C�Z���qǄ�����Ev@h7]Z�;�03)=f�M�v�G�8=;�X�����'n1�Hw@I~���%�w�Ƙ���IO�ק0mxgs,.�����`�]�Ȅ��U��_��������T|8�k��ݩ���b��绯\�Oh]O��k�:{�*E���5�W���~y�G�_����/M�sC	�K�_U
��NPT�d�c_��Gƶ45�4`Kz,�)^io��,��W���l
K��Ю��,�=FvC��M��I�q��}b
���L_�vD�tJ������R�_��M6'��ƒ�б(�J�/����S�)��;:���U���[����s֠v�c��
d��DOӂ�,� �K{�혎��k��+�kV�*�#\gX���>��Љ�t�On���h��?Y����:�e��x��p�*_���}x�gg�N]�i��r�ϽVȕA�P	��q�}=�;�g��D2�S��.<[ku�)�.1/�xK��LTO��E�-}��5Ҍ��$υfJƆ�8v.�C&%9 Q� Bn#\1�a��W�y���v$�p=VF�b4�H>�� [�7��F��:��q;'�?��y��H �5[g�U����H���L|̍K�\9�Y�J��2f.����nx|h�],n-޵~w�z��x�_Vf��Т��d�K�i%��Ֆ�P�r�E!�tV{�X��=�6R���<m��{Ýˆ�XH�=	�a}J�j��YB��/�TB�(|�)�B�f�9Fӹ�]�>f������^dppHV��pE]<х/�t���h!p�d���;���l;u�2�)B��l?�܂`l��aR��>.���W�|q����q�/�8r��O�KR]�1�ֲ�m!���bfCXR��Qե�seBo��\C��ki�l�v�nǣF��
�������D
g����2@��ݮt-���z̓�u�I�,�~���!9�S�@���A��h���%X:����߫�ί$�������14i������Ųc#� �-�bbx�.X>}�PH��!͘3�����/ڻ�L�@jg���6
��}�DM,�L��n1E�KHS�W,�=$��>\�#BV�?�F�\d����Ѓ/NL�	�%z����� �1"*3< d�JpA�t$$1A�-7�/�ⷋÀ����󧏙����Ń��;Do	!�O�B�`0�pQ+"KE�o��f%��DH#���yEQ~�߆�g�ŉ���l.jՃ٪�Y���`�_�Y�<�b/6.�=$�:�b��z��_t��#<\��{��.�H����e��jf�E����9�~y����wu��?��G��|�C*�Dנ��xz#�V�V�4l�.����� Z:a2>���ϽwNm*e�^#l>	֦�����"�72k��[�`�q5�v��'�ez!��{h��&=�mt+YY��D��?v4�
ը�s�Q�YD*����Y�tPL������p���P�����.�ݙWᙩ+����[���4_~�����F��c�]���>e|]��������������~�1=�,���H�\�x8z�%_�X��6�0�_�Mg��t�WKrk��v��8ă�#S��w1��n,�s�/Y:|B���~��IF��/F�^"2��p�1����u���j&�u�ӞK�`6�d�2�~����{5+�"[�q<�z���4��{�9&�ly��  �ϒ��u>ƚ�)�BJy��%�� h��řx����f,����
��Y����r�7}/e\�L�ͅ�p@aP#����#��=�G�)��ߞf�֞ ���E�����t���=�����?}����G��� �� ������^�ު�I�+k.�{!�;��Y��7n]%�ʢz��.�](y�@�Mg�Xߧ�æ��<[6����o�V�vzs?0��gL*f�&�.�C�u+d܉D=���kaJf�4�y������9|V�\f��C]�t���P����j� �
�}�X����Z�_�[U5��;�|_�6c��x1� ���ɨ	�Į5|�֋j���x8��Ue,7�5���ŕ0���G�z5o�>����-NK#�?��U���g\�
�9;���/��?���)w|P�'���f�e���V<[bACt��e�Cv��m�Er��ض��(��ϸ�?RJJ�W����A���?d|���|����(\�{��y�I�v�p�`Β���d�w��� ����dR�h��đ�M�0�8Ə�pt�K=��A���8����LP%:l!DN���A���_�U�0������"U2��w���)6љ\���|��AK&'���!��[W���3^��<�/*����)�PD�;K���K�67��bbb<�Mi�!8�ۄE��]v���[A%R%���ZGE�����霴�4J��?���DJ�d!�5��"@Q�X�!bO���<�f3�a(��P9
+=k����ѳE�T
U��
�����Y�|rlO�pW�6�|�	�@fG���6��[7�|���S�����F;�
���L=�&S)��������f:wR�$.j.�Xf⤘g5{=����$�1��)��+OBd/�ݾ��G4Ӈ�h)v�\����-�*嘏*��ӆ�,�Eq�,���]&kz�B�m`�9wNl
�x�f�KMeê]��SE$:P��,�)T巎5n��F7V��u��n�E���,�Ǝ9�.��'v���3�9�Y��l�p?�Y��3�.��[�������==�L+ԣl��VQKADE^��+���ܳ��O[d�v�Q��6�����[�-���i-���T�����E�RЄwƷ���i�����
	����		C���W.P	H�������&�'���0�M�BD��
�<q�uc��r,���"�f��ZJ$�F��F��l8���ABB~�.
��l��y7ۻ�H��x,��P,���)����f�S��o�����i��ΑV�J�+Z�^ ������>��Ǹ_N�qE���YoO��x�+M��ӫ���?�Ů�C��*QCW��1VJ��М�[u�o�d��(8k4[��P�-���lw%[�}�ޢ���Z%���djA)Os�\��8@�_��=m���踰��#xg����1��؟צ�3`��Nr%��(�v?]3�b.U�T������ޛB͞���x���N~m2^�c�[ۊ���Z Gl�o�L�l�v�F����;�.������D��*��9�DR���7Z��(����E���IR��D��c�7�-�r�E�����{\d�t���)K���eũ��N:/N�U�	��2��2�^t��_��cK�=����x̕0�"Zk���3-$��ȕ�J
 ��̳��s�ƍv�}$T�/��%[w�A�x�{���k��3h��Te�h��KDϨ9�-��֑6�G3c0��בF�Q�Y�i�`�#���>����FЀ�#��v�7��-�D�1c��� ���&s��c��(I���2��@ofY ׶�x6$8��.�b�]�X_ILk�:e�]G�m����oi{�����UiIfA�����N�$h{�Xw_׼\g�X�w�~���t�<ic΄2�uB���U���/�A��,�*{�SJ��}��|�
x@K����݀���4gD#�_�l�s�y�lr�g)4�F-v9��,����m'@��܇.(�׹��V��b�$���3��%�Y��EB �V?���4����¬������B�\fc˜��������m(4��枹����ݗlӂ*f�Ж��rrÚ��B�0f�`̒0��ռ��?�S�Q߫t�=c����F$��8��؎�<��8N��}�%���a�5��� Z��Ք��J_��ޛy�J�=uU�@LS�M��HXr����wԱW��p�T�s�v�E ��RS���X\D9�~B��"�������,�d�k�?AJ��Û2`2P�+�r���dq���y�'�3�WbV���=~�Q-�\���(��:r�JQ�P�H��aΓ �2j�P:FLZ�c� �����:.�pּd4�9��z�K~�o�D��/,����I�^�[e�U�'g9���o�.�R�-�]Fc��Y���x�
S�U`"�4��(Y�f[��Ǌm0E��ՒZe�Vu��_����jd�֝�J����ݞ���a=�E��ns�\�{͓�> ԁ�� ����A��?\&�"����y*�g-���UYR�'��p#����2��o~�/o�w\�#UE�L��=X�U���Ikɶ��p��	-����㝰��"�(r�r�Ee?��"�C��Df77��}���9Љ�Z���7�)	v��
�H�"�/�l8�of���xxy{�� ��e��FsS�܋�N�{i��
����8ц&j:f����g1��3ȳ]4�41��t��`t�� 6+`=�p;�oO�i��H�����?�����m;)���-�UBp�"�h�CX�{�uc�ɲ2t)���"������"/�s�6N�)�4�o�}UI4�D���+�._v�R��}�W @z����!t����ٝ���;�����r����X�R�*Ye~$GO�5�~WP�
-���Ny�J���������@i`�%̲S�Q�Ip��7�A�[�XM~�B���R����_]���j�8�ww�n�a���
�C�<��9j��Si_��sޗ��p;���'�ߝX����aI��&��K�p�I<B��P� �<�K2$�I@�L�k��F�?�}p�}��*�����2KQ�n},�|6qR\���E�GH��Wo�%}^���f11fZ�)mr�mR奵ٮ������ó��߿Q��r��`���~��I��s
�ҝ��Q�IG�t�ʆ�L~�-7��(H�0����s�B�y�Kh�ϴylO�Me�{'�ȴ�i��dk_���B�p���Sw{Ð/�����
A)�@
�CQcY�r��ٴOS����Ы{�OA=z(8J�~5k��xKP�ݗ*O�&�A��"1],3w�R�| �������&����FP�Pb��;H �����׸��Xn���.�Wg>C�yY��{�c�Mw��J��]V�Y�@��������p�$�J��=وF==aOI�H���n���3-Ms2$�&�Ip{c)C��~�N�c;�|�x��ٜ�Dx��&L	9x�po[T����}VK�ʐܸ)�y�B���ӓ�aF���{ƇA��;Q%G|$JAf�ÀR);�KY*,�db�!mJ~Ә�P@Ҕ�B�����ɉp�<h	:���b���M���~o��b먘2�_��>�V$�!{C��@����I���^gf�_��+%a�� ��{�T�)G���A�\�2������ É9A� �S�!���Eu�7f��:�<���F�G�1]Ǫ�F;7WoP��l6ۅ���y���؝�#����_:� KY�����񺗙�b]��վn[x3�V4��B!���]��&*V~�]L�ȕi�$�Ls�|�	�"��ɠ�T�\��_�Yf����.[���l����$�4)]6{�Jͧ%�Ֆ����\�}T]����[��6�[!KɎMNM!Î %�.\�c��C_U���ڿ�X	2o�V��e|�i��Y��h�����E��BV��p� oN��΍,���^� �ɨ���:���ܟ
��O��b��A�碇�		�ܲ�Hb��{��Lټ��U ����I<����Y����m�?<3Dc?�)dy�i�i�����wG����F"�ܤe���X$��8v�a^=���My`�r竢#.�.g����O���3 p&C��,���{�qd7^�Po@��x�L�c:o	�!�Vk�޸��#gr2���6��W��� ���\�fS�� J��$���-Xc�-b��IV���y�/�񤳝ߎ�+>^I���4���q�_����:����V�#�s�\8����k�� a*+�jċ5�,\�n�Cu�;�xkõG��:�"^����5�'��7e.�tIC^Ğ6c97�J�4ʆO|�>�D 4fB-�Y^�0�3c�	:ne��$I*G�C����uğ��D��-���hR3��I��.k�֌��v��_|ʖ"DB���E![Zш���2� �������E�@��&�v2N^�$�"Ӕ�4)��f֘�fp�w:��J%//�����"��Yy]?����a-��C�[����}Yau�[J0I�����O��I+v�|[m$AsIZ,��¨V.������./ޏk�at��MRR�A�n<��8�h�5��;��Rg����?y��2��ܦ�ҕvdPh aq�KM�'��i�g��~���v�Bח0e��_��������:^G%m��4Y��콓��>{���g67Km^��#����P (6C+��6���x&e��%	�b���iX@�^7J��M�No��M�V���D���q(�Zi$$$_%>����ï� b��wB�_1wbFT./幗��^O��º��Md�K{�C�Edu���/ӠI�ؒb4��_��)hiF:��`�C�e�s�<����h�Uc"���ل�F�''Ypm)K.��a�zۭ�7Nq�;����#�\�FmH�v����[Fj�0�e9:3#�����gQ��",׽�e8��.2s�VM:t�s$�:���_��oj>�C+ 0�6N@�|iH��H,׌�O�����'�0`���Z�0������/<ߓ�;����{:���k��e�������8���T����JV:-��aTJ.d�3:��c`)�S	�U�IIB�W΢F��oQ~�;����4�'��U��4��F���$9��uW�,l.��)��^(&�@xD,N�(���,+?(z����d��(D��џx.Q��9���_Y�}!���u������3/7��u6h@�����7��P�(I����ڄ'�H$3e�\���2�'JՕI�JM�C���W���Y95�Ǡ��Q��k����+�W�Y��/)�<��L]�V7�R�.�{��f��v�tZ7������&�5�q[��ʫ37�f��~�����*��v�;'�}���/��I!/[4g����	AܚhCN���[>*�V�H��A��ёb^o\y�J��⽕�D2{Ռj�M�i�{7{y7oPo�ƅD�C�;�$Ii�`o��0(��F@tww�!�A1c���Z�t��P
�-q���D�㊲�������ǽƙ 䠹zE�i���Vv�
�)]��=�L�_��L�M��"�	sψ`�ΰ�;Ե'=H4~�K���N�ьu��+�
<��x��3u��A��'_��>c���o0
vFJe-^�����8<m���*V��@�N��(�O�Y�������9�yW^eI����������2(������N���� xp���Np� �/��n!�����G�����۪��;gN�s�{:�J�)i���/�Tf+ۊ�F��_�x��^�6�#;".N�FB���a�W��P�w;Y��~�w
��A�shf�Q]��H�8V�}[�?a���Ȕ-O�׍u�--R^x%�"�4t��dC�=G��T2��?�7�">�V?��Q�m���W��9촄f�P���¼u�=��h�z��>Y��q��,� ��[ͷq���m���?��$�tdM���f-lUv2���ݡ��
�}�v���@���D.^2�$\phN� ���B<?@�ٳ-Ļ�o]��,s�P�ܫ1��$����v��c�]���"}j5����?S񦄳������R���ˈ����N�����'7`M������_��O�~͡��jr��E�
\�������B�jJ��X`����VK�V&��*� �$�3������ڟΛl6P+u��|[y&;5���؃ҞG��z�6�F���r��h�U��jdF�z�,)C.uRLϡ���ȻyGt���?�5�Vg���Ǽ�vk�?��������-3#�J��t��ߣY�Q�Ϫ��̘T�!�w�QFUO`OG��D�W��/>p���q���b9y<��=#Q.��ƌ��r�1 i,5��4�{3���}O~��y�y||��Af�g��WT+�
�Q�S���*��"Rݎ�TG����J��d��)j��P�_|)�k���:�TR�����t4M��Ea`��5(ͨO%;���	�C7}��
١)�0� 8{;�N�~����S�!
�2�t"^�9������5��VIg�w"�b�~�7�O����ꎿLG�>�?��٧_7tѻg�q��J3g����,5�q^^��n����#9��iV�k�d��b���پ�(�����%��H�� ������r�B��`��c����ӻ	��?l�"G�f~�Y�\>R���o�7���'?B��x���wFҴ�4F�C�q�G��[�( #!�hX�!,�X��dfh�D�C@f@;o�\�Ia��@��g��0�@���{�_D���~���1��hj�����lZU��kv�o�7O�ve#�So�8ӹF~��]1�j_�� B&L�	��i�G*��]���L���Fl�X�=�h�kQ�M���P)�
(P��C�3"�/~_�C��][Mv�W�0ߥќ~t�f����{$���o�����.N�޺�ڵ�#��?�[6�����2��o�C5�|��G.7��#g|0�j���|9�߫���U��eXl3%��ZW��UE)�{��!�a�� �����c���� �-�P��T�1%c�.��B� ��M秐�zHE�-T���3��u�ۍ��Td�\���D�b	K�COOρ���,?��8~=�3���ӆL_N6^�:�2�y���ѢD9l���5�},9FnYԱz��k"�i2��{k56��@#w�Ä�Os"y�D �6g��z���"*���i4�
l��䛙���\D����)�*� '�`������O��@��`x.y�D	� Y)V�<�g��|5�<')���/���\�H�S��?��~],N��tV���W�	�Ӛ:Nn�{���~+jH�o������?���菰c☌��i���Ή|�*%ַ%�H����a8��p,�'o��2��w��G�O�o�9�Hm!�TŒD���]3.�8e��1�i鼵r��6� #�n�,ڹ�̗8�]i��$�/̀�B.�3�� ���É'=�o�������v��͕��[�_8߫��4Qr��`k� ���$&�u��� ��]�b��! �d	/,G�k�߬l���� k�j�Յ�-����I~��'A����1��u�	7'0n[�#��1����E�SX��˄�-�H������FF"�]�U�<�������0F��ڢk�����^Qyp��<����;�`��ف��kJ�+�#$��눇Ҙe�QW%�
U��i�5Z#N�����3j'��,�m��f��ʁB(���~��>_\$�<��-PO���ɒ�=��*ZT��۶_��`�m�k��� �(� מ��V�S���,L��'�; [B)P� �!]`�E�����f�(��~G�]�NU$CѤmr�-hl�A��0�W/��w7ǲ'MS&q��k]:����m��)I$�[}��K��t^�o��s��g����@f�u�MI�م+���G�U�-��
�Yh�w����ZDڅpR�j�i�k�q)^B�p�An�RVG�w#��G�n� �[/�� +"���<�7���I_��Wл+.�Z��\�涔�������C�Y��Ĭi4W���_#_�"P%��������(����ƺ��M�j7ң0����dG�Hz�g��lRoC����|c�rjs!$�S6ՇƁJ`�ۅ��������L��v ]�մ��>7��ؔ�FNz>��IwlV���[u��2�G�Qff�����Ν��h�T�Z��&����А��鉓�#N����ד��'U1���)F'A�J��r���"�/�����E�����GG�v ]
���GV�Q�iLO��_��)�o"2O��cV�����5�{��k�=���={��R���U�O���F��ǴХd	q�t}x���X0.c�3�
X�����%�U�ǚ&�?Z3e��d��5O%�����w����M���!B�T������*[�~��vŜr�\=��e��@��\h�A��Z�~J	��HQ�q��������Ε��/~������;���%=7�A�a�Q *X��mrn�;}�5�PgA���yo<՚`�Gz,Ot[؅X~���X�� �0U�<���tujqW>[k|�����`��ie�ԔJ�k��=KǺ��/�7�^J�sc����K�L�ZLҋ�r�d����׫jM���r@����4U�K�nOZ�#�q*�+$�	�JR�|�/�(X�����_w�uh�mءT��0�;��*�����������H!7-�Ӌ�O�� 6!�o=�m.��Z;W�_�T�Y��`Q���y[����%�_�6f5�8��%ޣE��7�����2+.2w�N{~0s��.���]Aɂه���&POR�����V�˩��U�5E��$=i�%�m+ jEGn� ���"�\��ˀN��s��<ƣ�Cξ q��<.��<6C�/HS:�c�^��S�_�;RO_�����P�������R>{�/_0����/'B��Ҩ��*n��V�+����n&o4yH!CdQ�Q+�"�l"�i�)٭9#T�� Wd2�r�OkG\�f���+f�ƀh?L1�ƲYG�zOn�7�W�Y�����_5!�CUD�X\kr����ح�l*�I��=��b�(T#����}Gf�!���g�@*<2S���(h4��zA��#��KEH���j��8tO�'��(��a����E�Zn/F**���Q��5�;[h�ɧ���v,lêiҪ)�Y+�K1O9��Q=�*�q��2�w��i%�=~�?D?�"-�q�c�9���DH}�.���( �����=��<�75��8,KÈ�Z�;	g����<����&��c7 e���ؿ>p���x �v��	?�n�u�%Y\(�r�4S��g��i���
���sz5.�Y�������B�=�W�3�G����\�.���f�)����4��0�{2����P�I�Ƃ���Q�_��I񩮎sD��T��dŜdÒx�U����%K#[[4VRHkZ�,�aV������)Ki:�j��X��%,��b�4ۜU褦(}҄N^�T�a�6��i�����o����������n*v<���AqR�����v�;O���@����矿-{KJ�<�G���Q���m̿�����]'c	vH���,~AC��$00���V�V	���E܇8bʫ!Pl>�W�������I�$�@2��ԡ�2Ǆ+���NXNQ�`�^;���Q/����ה�1�`A�ғ����YB��E�$�ϯ�a��^nLg��D@��=�uEo�:qĿ��^�g�:_��dg�UXDr��(C�(r�y��ZJD_@jr���L+.Ӈ9t�r��c,�y���(�r4戀׾��� Z�B(G��c��S [�6P8����TP�	����f�v�A��Q����i�T���JA_?�,�z8i�*���=P|�� R��ζ;?�����#���J� ��Z��嵎��N�S��;@|C\j"#����R��T���~��A�����`9���3�aROZ^5B1�)�x��;a�?)��'��m׼�܇�|�X<��F�a�6��H�zX����X��z���������S�&X�"���y\��A$q�����Z��|�O�l�yР�V��O���r�ݧ#!$�r��y!��ÙG���0WJI#K>;�*��/x�,#7N�>)��c����jo,�,�y����ֈ�V��������D�@+�Z�ۼ�b�.��<�z���:qJ�fc���X�,��Bm��R�6ÍA	鰤�{>�pZ�װ�ܔD�"s�T/�3"�M�|�f#2m��V���'�M�T��Zw�&�(RN�X)�̡-���g���C�}	dVJ4H���΂l�T ���^-,^UU�:U�Y��kQ�����^g��{C�k?���~kN�+�'�Pg����进��	��=��Ԛ c�	m�ʧr����isO�t��*�tgEn���m!I����`gM3�CuX��f�������y�)#䲈K�r���`4����HN!�w�d;��(rt��t��9F�P
ۺ)]Kۑ	e���{(��|�9a�"�Uʌ�~J~|�T���<���X�l�/*���:��m<�O�ȸ0L�.��ʥ�~�)0	��Z��;`�ӯv���~>IJh}��Kc�7�z�zx;>B��C{�v�V�����������3q����"�iK���`�x�?�����G�i�~vX�Ȭ�k���ؙ��tW�܉�D�/-*���h(q=*�fϜ:Գ5 _[��:_G:�Q��_=}��6��ym��4�v�!� �� \.�dL�Rw�&�(�WC�&J¢�S����:"�+��'&t�v�P�H�X��ҟ�n�"�2ic�m��h�Q�8Ԋ�N����sdФBY+�#��T��^0��.<��6d,�G�&NO\����V��nR@((N���:B�1"��&���DȻ����$n��W���A��e@L�\�jng����U�	���},t;!��0rb������p�;��mW������ǊL~J[�k��Q1�"�a�j! �[���0X�cd�6v�r';�!���nsq��c���Zy��z�X�#��UNf�7���)�l�V�!�s��� ��$�v��ST>_A�՟UE��Q���WF�������.��)ݒ�C������/ٯ�N���e_|Qtٗ������oyl��	�ʹ-.�E��Ն�پ�̆�-kn���E�T��B�,+�d�H�ȉS�i��V��V���8��R�D>G�|�L�L��MG�I5���0n��Ã'�UA�p:60ۋ�|b��˷�5�5��A�h
�B1�M�b��Ul�L��O�$�bi��C�X�\������oMm+Z���&(��ϛy�р���\��#�!nmц�Έ1^C*?n�u��P>��$�70w����jE,�h��>�3��(_/Sn>��n�%�'U��L7R�RV~�;���<�,���an������ȣ[�����]�dZ���G�uيI��H����h��$�}dNX�ny��Tst���H[k��vBS)��U��W�R <��7�,
��h"<w�,۴J>R�\(\C2.�2`�a��Ͳ���� K�������Béi�O|0]ք3Ě���\Q���o5Ormk;�/ng�Ѧ1޷ǜ(�:�V�
�a���U���hafMRvdZ�F��[´]Y���$�����ÆB0��D\w�ۻ���3�ݐfiJ�Ls�r��8���9�`�p��K��9缾p 	�
@9@Ҥbx&9,I?qc����)��ykiDE�	��X����DP}��4*��������F� 5�L��f�`��*8 ,�AP�l�S�����Z���[�.��Ð��X��w��?[u�G����a>LM�9���\�?�-M�ܭn_�r�<�>û�,�vt����ɥ�P�n	0���P�|g�vEXY���J���6�۲-����B����h	
	c��"�0		��U��/�a�8!�V�P�mJ\)��ѡ�d �l�WC���t?�R��dzz��3���p1�-������+ fD&�p�F��:L)�*�,p{?����j�c$�k�'>���:�_�g~��%����G��9��ȟ��E/��01�'����fa�9�z�y���.A�g�Y�i��>䋘<.M�����w���eX��7�w��!�>A?}&�[~���1e��f�����TP~������|�ML��c��ȳ'����2�G6W�����	��U.S���t6���ܳXVWv�������]��z�1���������t(N�!@
/SEv�>�){������ƀ�֚���?�.C7�.$u��;�x��Fì�<�O֯Z?i� sXnD�@���<��q]�z�������T8�j���u%d��-�pid��"6���v,�����
�a���!��z���u���*�W}�m1��f~��������YT�K�i~&�@���ߺ�N|P�(ʗ
��)���qa7/1��IJ��+���G��� T�CXLVa�þ��O�1�w���u�/���P/��c����2?x�ķ���%v��z��ۯ���'��_��H����
��)��D������	e(Weï��q�()�=
����%غ8_�g�,�<�^Т3�#$|E?e놵\Q���&�w? ��7~כ�Ԧ��
�/�֢.�i,\��Uu�>���5��e�� R�[�vF��v-+� �WAK�赀:F,M��Ӆ�,S'���	��G{*�2���=8 W��")��	13��o�t�guU[��h4���b����n�ɦ�n����i��:�V����Fƈ��b��7���Fg�ے�O?J�(��_a�Ϝ����

JՙDQL��g{�͙�Th�S-O���޹������4�� �2���G,���	Y3	���V$�<�
�	�㣩=Cc�� ��)��_(O�Z��f�[��t���Űu��8�.rbEe��ª�e�<c�ӳ��?о�[�7L	�9��d&����@#ޝ_����I.��H��:
#]*�>�F�j؜�� �� r�P ĭ��>�+��ㆉ�4�l`�M6٬��Y^I�	)�L'X��t������'�_\�H
�J���k�Õ<�FxX���,^��?�+����V�`�&��%�|J7��.[o�D3����M:F
�F�L�9	�@�*s�Ӑ��s���VŇ�m@6F�b.n�H���u�M�"���~<�](��}B�탛��nۿ��&���8�S?���o�ylu8m��a�L�+�%��8nq��w�F-�n�Nw/�,3�5�9�b��U.���HI��A\�7wh��<�%��$�T�'O�H�{���#�3=�D�9���W���)o�2u&���S���b�S�$�0#�Ɓ�9r\�Ō����X�a���; ��V�F����"ʰ�O��8�a���T�iJ�@�<�L�Ůp��?N~�����~m�j�G
�Qێ"c���5���1����z��	~���oOC�N���3��)*����缫�0�V6+�5N�z��i�-zf!@��}	�L��ό3��;��߇4�W����u��'�)���?�idMr��:�(�&�t/0����#E��3�;5��՝s��'�B6�x�'�"H��◲���\):�����B]�5��X?R�!ԭ!�e\ ���~��j�S���H���R���
ϩ���>���t�\?B���P5����?G�w҂�L��O��-+�r�+��1hDX	�P��N��������W�d1R*��h�0������#�k�g4QM����8��+<���4+v)�kI������\ݨ'*8�&����1���ۥK����f�Wr���p��1���őV��F97�SB-�K����E�2Ɓ�9�G���m�g�_M�<zH�ṙ�!���b`
��h'�Re�?v�8  �Xf���8�$��B���c�W��?
�X���Lo-���87ɮ�{��qR�2��+��9�q*���\�v�y-ivɬ�J��ܼ����+��Y�x�c��Vz!YD֌��#1�sG���o�~�/^�$��Vs ;�&�U:0����~�ͼ�j1$�վ��[�2T�a�wW�ߎ�l���n��H���|���M�1KV�[��`/�D�P� �o�-�m�؎��a� �'�[�;͌M�m�H��"eT�7�������ʞ�ÖO�y�/ ����i;����Xl�3��V�H"��hι/�X\v֭���Ko�6��.�X>W��U\,[Yܲ1}~�_'G닰�>n���[6$M@נ�Fݺ�9
ПI�E�4��>[�����u|��[W�^��R6�����>�l�����q���K��Q�Q!��u�N+�3����Ay���ˆ��0��
XmI�B�`3�im3���]���[>� �77h���k�|@��RGn�FA�s}��J/ C&�j9�a�����1��=�Msv�5�JpK4�}��&���`�ZZb��:��rE�e{�����V��I�uP�'�+��1N���Kd��G3�^��}:G+�K�`QD�/h�<LDDmt˭Y����q�G8u��؋�}�?�G���	��:��޵��3���"_�2��}%Bi��$6x�J(y}�z��Sy�4|�2�*����/�f�M?;��2X��[��r�� �^ 0�w�)���tH@~o钅�߿I��wځOMڡ��#8�9���'WJ�I��]a��j��8*bCO�%is���z�
�v{��h6%Z��,P\#y�i_�ӫs��̳k� -��Mm����MXrQx�ob1��>ih��r���kJ�x>�.��Z��z0 �����h\ڡ�������GLX����bJǵ9FnK�D��^�Hl*�S��DI�Gi&�'�\]К�ЮКj5��O�����j�� �Xj�����n*Ȋ��
����ǖ�d))�$%p��%����A]��j2	�6�?����(�FF�<R�yBi�����ƫK�y�Q,s��F��N����-7f6ذ���~#x]H�Pft{J,����&:��i�Y��@��Ϭ��բ�e�b�R�n6��.ە���/�o̎��߸"7�~�*x�g�"XT7��0��-=V<�m�e�{�r� �.���"����y�J$�D���6�k�1�g�M6�˖2é�f��4v�7u���Mȝ��[�~R4�*��-�C��/��K��9�6�l��c�>9vNԭA�Yz11���%Js߄E�7�^���~TFa�����.J������i%1|�"<�R����ؓ��q'K�f�1D_���wo�Mt��/��NE��:�[7�4����/E%�Q������S��Z�ąj�E+�	�IJS㦑 
("%T��-J3�٨�i�y����9���y���������u�X!U���E�`�  �jr|�2��lZk��=�f� �JL��E!�{ɗ�q����tl
A�){\�%Ri�^|�4�'V�|XEq9��\I^��ѻo7���"�?g�k'Nݣ���y�iF���,{��R�ۿ�u�3��Wb����5l�4U����Z�Q�ğTӘ����4�Z���W?@���*���/�Ll&C�E�NEU�K����bV��nX�1SC:-����Y"��£n�qV0n�h6��/�!+��XV�I����9�f�x?��NB�W���E����?^>!��~�B4���ר2b�3O�L����vS�|�6�v���w���k-�u����������%��\~X��Ԛl��=6{t�&��w/��wwT���v��b�4�@����/o1�w�.V��Y�2L�~H9�q�8��I�E$Fx�r�����9g�)O�+Q�)O{irȓ�4�Ŭ���X�_�4��ċ.�I�L�,UZ
��)�gv](}�ip,i��>D۫ʕ�]'�]	��\0�* kD2QF�?!�kߏ������C���=�����i��:s�C���ĉ9&70��OL�Kb���u��v:��(ɬ}P+��O4�7vPi�y;搏G�2b������9>���au/QI�B����nk��d�/�ԇU�i��09�f��4MeO�N�޼%({ݕ��4�6�`�<<d� #�U�;�+?�ֹ���e�Mb�;)��F@^�Bw'm�0<���7yy[�,sҼ�7���=��b�Q�AG���`o��ǢM��?�Kz�i��r�;ݸE�G�i-U����.B��=��\���+N7sRZ�o�d3�~��B���/cڄ�nhb�[o�Ù=��P�礩��7^�sZQ������	������Ǿ�+���l�U�Y��0T�u����-�\&V4*i��̝6��;RK���.P~�l~�Ŗ���gfm��۪ ���6nQ�[�Ap����k�ht5���	��~��Y��iB�om1�w#�^�A�`5�+�7���D̊����?t��1(��8��~��G��ݛ�T��J�$H���k�y��+#����o�Ո�ۮ��b�:mr0K<�*��MI]�A��"�8�y>{�zC����SX�˿*i�l�g��������ZҎ��cA����(�AL��`2�b�n��^+��4�E�Y�,H,>U��K&aj3�.��W9���e��"�B��H�f̝3>�]��g9���kɛ�/�-e]�^��D�n�(� crp���1������L�,�O/��qz�Mپ�]��^I���~�cF�����!ֿ�!������ӧ������F�$���Z�D�t+e�=;:9��C˙?4}�rHj��<��u(���)� N��Z��4*���d���0���۲5z�R�_gs������w����ha����nI�Ir�!X�L�2�M�s�h��RHPhG���ᧂ%U��1�4$���iH��Ӱ��N������P�����_D��m���
c�'vs�wco��*��0 %osC*���f��A�I���2f�@�⼦����J"�؅��������^�,��ld���2e��߶���ば�:���ט��*DT��}�R�qŮQ��ԑ�P�H�S��@�
����Q"�����䄷@ e��l+f��+q�0�����e-��;����s�}�y{�"���� ��҃P�-���r�L������O����|P|��.��~ �g�Fz�|��3E�rJ��R��b�-�ȿ��%���T�����]d0�X���Z/!Ȼ���f�!R�l��,* ��#g���p���3z�u�����Q�dK3m4^8b�w����
�x�YZn�8�_���]��k`G����QX�R��|�E��_)��9ۦ�]� %M���)���b�M���������j�8cD� ,'7�4�}~��4ʿ�z���_g�V�;�8��	 ~��h�\����f�Z[)5#���"4)��������F
T�ʙ�JM�ۀ�հ��t��>=(Tf�M��ۆ�nmp�6�ٜ��ܪ��{��=����{����B�Uv�lv�-$�T5W�C�y��Y
��C���Q�V�ߍ�Cl�H�]��gƻ��
��k�n/A��4!3��.'君�oi�����M�U�AT�0����y���6���PW̃��a#����xnQ����j)s��_�u��g�w!�v���/� =�R3�N��Ƈ�`��O���f�rLH�W&���W_�#?�G)	 F��P� ��V�u��w�5L����8�,�v'� 	��nVO2��o��ž	���׿��|m5�|z�2U�综�����,6��K�̝�S$� nj�FMM]�N��<FGM�φS;ُj�/�Pu]C!:i=��[���Ŋ���^zxXb����b���HH�-<�FM�A�+wi�����3CN�����+�������J��Ql+K���~�<��sx��3'���h<���|Ϛ9_�y�[���'d�$���j���zÆp2�3E�@q�t�;M���p�hT3�������Is��z$�׎�Nɋ���*#��*�U$C�����I�*ƫ}O#���fq`�fi�m�����e5��T�{ho���ŷ�V��"���b?�p���)�V��w����S�U��,��y�����M&�(���~J��X�TI^�b�?�����$ �|����ϲ8�N��N�;y�4d�E)ډ̴@AHL�����r�Y�-�r��@�v�߼)(f��es9"5�t��=]/�-/]iM��g���ׯ=��������4�������w!�h�/.�D#�T%cGٹ��k�D��/��g��oB0kT�L����Us\�k�,��.��_�i@%��v��۞8�� ɤA�F%�p�?�/�p������M!+BDD `Li2����e/PtS��k��y��L�����F�x�����'n�8gx�Ge٢�C	��[}+�m+�M?���c�a�ܼJ���mys%�����S@�� wg蜟ĭv���!Aң|�e9�ʛ��f������������DVT}�f�]�4��Ec�=0��]���Ǵ�~�?�v�ɺ:6�T\��5�Y����%0�[6	9�l?�3�Y�ǅe����](=�r�\���Le.���?K�h�Z-(���f_�A$�X[�J�c4��q�u�)9_���x��K���iȌ��xnLRntЭru���*�����]貔N;hge��L��\��TӘ�\� �<�H��w���'-�ab+fi�'i����D3�Q���e����6� ��{=U���U�:�����)T9E�(]/��^��Xx�m��̕ S�eip���>5����N,�S���U
�::�M�fũZѩ�>�	�j�M����!�6-:�����q�d^�x@{U���O(C7>P�O��;�](u�+�>�qo�Ww�r*z}�{�x�p�Vw��f����o_�{��]B,ar=���գ�K+�[j���+�BO�ǩOZ�ӯ�}ܮ4��>~�
��3���S��
� �D��"��M�!˺��*LP?б�x1o5�>�ѐ-�|��I���,7-�\	�; ��S�z�]��K.	�������9�K�m9��b��(V�CB?]-��rhg�x���J����'��w�Nb??��
�N��d��^B�TQ�߲G�f����M�֭ݺ0��4���R�5�*�����n���[uG�huS�l_\�X���Xȍ�-�[���R*��(����0��·���I�!�:���];;�Q#

F&&0��2�)� 1�ؙ�/�;C����u�a��ٴ%��t����it�Do�:3>#\�uF���Wk��������vn�n�-�j���&h�7{�]l^��&ƿ���u�v�i]���6�j��d���#��7<���s���
�<:�� \�3F��c}X�j�Pj��.��^��(y�ˊ��>���_
G|�a,2Bl���ih撝��9QB�H�s�\�rT%�0E�j�Zى<;$�|+Xtp��]�V�����1�  {�����Mk��dnv�B�_їB�+�W��Ğ��$��4��$��[���G�Qi�7����?�0nf��w���:���sK^-"'P�Va;�Rp1�U}��uM#N�]1��q���,�|!��sKؽ�cwB����|���e�'��D_d:',�����%I|����e���ׯ+2�����4��(��,��_��}C+�v@@����\�v�ڐ���~��Y��I�k�.��Ҽ���M�YK'��z��㗔�e�Vb�^/b�Q�.&e`]\J�R|� �k��Tc�Kq}���q����%eh	S��\����?���wL��rUuI5���Q��+Q	>�/�c>wc�/>�^fK��[�$a����r��F|��m"^�SY�Ci{��/�7JHm�G4/'��k�!��וk\M#<W߸��[f��̒D+�V�Il.�x33ܠs��G�_����}��I�y�ta�}[��ƴ��Y%!`���} ��S<_q8��	3�6|�V�"�F��qs'�o7�S4Q-�eHFo�j+la\�8�&�%��E�����l�)�uQ|�[R:O�,]wI�C_��ׯ"�5�A�ġGŎ�s�flM�g��2Z?��R 1��u~ѿy��[�v�`L�b'�6��q�Ww����O�7)���8����y'A���'�W �F���zGM�U�J-MUţ��W��m�&l,t����o�6���_�}I�E�?tD�,��։��k����嶐��h��N�) ?Od�����b����oy	��9��~��'aX���P��ӚX���}�� F������%���CI��n�*咽���CQ�{Q�3������̜N���TP��j�lc���eA��GO��o���/��P���ޮ}�0�>N��YB�oGՑ����������cq�S�u����l����1����La��2X�Q�8r<�dyR��$� {6��
�����0y��M�!��K:
��=o��T����	��An>C��Q���s�Jbᠪ����:$�w���~���%(b;GC��ƜF<*�p�w��'���G���:�?fy��ۦk���ɫ�N���ț:q	�,4<\
�]����E��M�[w[���Z̷-;e\��\�0� �s'���1���Ҝ��r�� �6����r&>n��쇱�J9�<	�%�ݢ��>ٵKQr��/K�1���������L��M��J�+�b��	DT�P�&>߭X�С5k���R ͈�}.e�&ٸ%m�ޗ�����q��Ք>�R���w���AC��#(�͚P=l�D���{���N�6i��_u�;$Ia~�Z��W]k�������6,V�ǥ4�z(R�����H���8}o)[��G��C�:��)丯�#�~l�|��&�(Z�k�bEIQ��l=�o�wKp7�� e�H��K�s��H�H= )MT�J����.e�N>����U�;j�!	>�4P����4�����-cz�9z 0�"�:���C ���~�2��Hd2A���Ug�W`״�V
_�� 8��;X'�,���x�x�.	�|���?�4$��k�����] 	�����&۪i�<�������uNO8X��5>00���8��ַ@e����N�L1�H'��Sv�����oTvY�v��Vq-�D]׳x�Y�Q�� �f��<�穰ء��h�`6�`�[�l��U�4�Z��b��P7R���pS�/�Y��U���M'-A�\�H�]A�A}zْ�n='Hۺ���ğ��7�3����H���d�,��¦���ȷ�V�*"5�˃˹��O����ƛ_&��WDl�*W��a8��0�N(���l�MF�_�xR�*�v�U�__�m�ǸQk�Z�)F�\�{��˲��(���x�M�}��k��e1�T�<)t҈j�]2�б[8?� �H
J����$����}`�c$f��!�{g2�	�i���DIf�¥�o6��u��`Lm7�<Q��
UdX�2����؋����`QL�1�z��>������2�Rqi�H��u\���֍x�Qㅟ@�'cg��1�,�o�7l�t���V�S؅�͈8Z�;�gp�Ƞ��ZÆ)2��2��!���ߒ������8炀��9L�4��BkL�����>��j�37n�奸LX�:n�y�z[��mw��4�֑�0�M��ր��� i�=n(�f��`/����� ,��i��Ӯ����[��-�=p��k4�d�x��c>.#<U��>K�=�k��N�a��tי8>�{�.L���G������G���� ���օw���:��5�;��w�	��ww���������=�꿷nݩ�����^�V�^�yf���}�b6Y���!M�v��S�S���v��gY(�����D*B��Y��mbp�#뭪��4��n���)/�򗵅����I�)�(*CE�����VbƆ�o$Gޑ7�6�W��$�#H�o��nY�m�1w=X7;���u�ܐOw�&8Cl��i�����?Ĵda�ੀ��pC��/�j�/DtGrtȻbēs2DN]\�j8%�����9����4K0\UYi`��`��>��OK��PyK�%�OMM��(� ��&�;!Ǖfo�mZ�m.���5WQ�3�|r������-���,�6*�@��߰au]���Uj7�~.����J O�uưa�N�7��G` U?؞�.��fy��1z�\�33!������hƲ���[�]'�}�2�gWu�ukED%�~4<A��A켡����*y������r]ڡ];3%X]�_qW3�Q�Xc�q�ud+g]�����I#�M#�� 1��������lb��+�\ƷV�jyfe�r\9[Q�y=β����]E��>C�v��GmK䍎�ϵ��d��t�-`k����u�m�E�.�Y��?guUƳ]��na8,"
xA|V�co���-����Ȉ��ͷM�ڳ	�̳0x;m��n}! d�p��h���N/{6Ͻ��ݝHTr�Ы�Cr�
UJ&�g"�γnpJ�t#$!W��Y�dd�O��kе�uYk��|aY}����͓鞇m��pP����jr `aa�x}��e��Br��Ѽ֒�D@��*Z��з��='��f-	���x!�����X���klR�)a`}kXTjl�DhƸ�9!m\�"0�6ע	�Lp��u��6<<��;0� ,h��`��7��([���f{7�W�R��r���͂��D��}���+��kXjm�+Rr��1����"R9�M�\��BK���?_���A[��`�)�Z����`�W2�0|��qĈ����3F����0?W�rA��h�J��{��LJ�E�,�#ٶ���N�u$�&�j��tm
��ܝ��n�7�+�·�O��е���Dd)x�D����,G�VS$��d̸	!�0�,LZF�n��2�?/pk�ԅ�Z�������GtU��jfJ&f�ʚ�*�H�r��T����9���x�>̢�Y)?�*�k�����, b:�Gw�-�&(,F>�p#�A���)��p*�����p^S���j��-��&ͭ3�`������ =U�ú1�.v�8�@��^�N�s��o����S��z��#�}�݊�iǗ�w[�oF�3��*&c�(f�*ͼ����љ�B�k6KJ4���x�ݣ_�޵W>E,�;���kd�7A��T��<�+���sJ�Վ���p�"�?�{6��ھ�~�bH9�O)a�`a�h�&�:���:t#r骉���LO��TE�v��v-��v�m֡ХJ�]w���"P_��� ;�A���|��1�-\x�~�R�+��j$5�A�#���}W��T��g��]R�s�P����w��Ʌes�1?��܃��_c~�/m��g_��o�?�{�j-1�S�ل�V�9,jP�9��`dާͮ�;�F�-����}�0�����9q���^�st�Ԑg��,ERAb�j�����q�/>���U��P���>$�B�{�kAp�D���p���u��#���G�ܓ����s߫�����gA��'��p;��
�*K7�����.��.'L�X�Z$
j{[��^7/q�4	a�u_��k��5�b��O0~���N���z���<nL��W�0������)ř덛��d3�$I��^�}V�ԫ�ɥ�Z�u�z�.�{���ѵD�7���D�dFƠ�'��������t����6��z)=��1H f�2��D�����\vϭ�үz�:o_b�k�������xY��zOY��[u�Wn�~�K� ���^�pV6�P���JX<�P���<�Y�P,_^�V͠ N�l����
I]���Wv��ڢq�M24@ @`�ӽ�G�;�{�i+~��>���;	ݽ�d�uj<�L֔ޞ��(�ˏ�:w=g5��b��t���L�&CL�����Ϋ�3��?'��u���ȴ���2܍B�
��#;U�%P�p���i!(�-�������D��y}s�>Mn�X��,$�\�gf�CLII�O�;�V׼קd%Cc��ul�_J�ϭ��b/��O圮�DZ�U��S�%���&�~�HSsdEB��M��Z�گ$HU�:��%�e�{mQ�P��'\���x���c ����b��L�P�q7S�h��=O�� ��̀��龥����Z��$`�V�A�w��c��j;�����{��{O打�[���Q ,�ګ�p��Qf���Bx�G���D8��D��dw�ݧ��E𗑁��M�6ү�r�ǈ���"}RA�dr��uOO�����}A�����*��F��u.��*��O��/;+��ý��U�����+՜�hx
qkO���̸��Gߚp���V�P)��3	T�S������	��s���&��S��֭8'���$
0[�N�)S�7 e�)��d�_��ן����a�[Yv5}�}���$a�$�C5Gr���g�'Q7	J��$R@V9�U>Q������U�k���{O��5s�L5/�W����~�~������De��q���7��Vag!��D��⤕��@{�Vt�>D���(��}�=�߿�ds�ge��<�N��9��Z���f���
͸ �V�fX�X��a�!��_�R�M��4u2~��K"t�#��Q�T�ю�?�RM�YN�=�(��-�W]��34�)f:o�ʦ�͹k�˥� )�+�2�r󨴲�,N(��sbVM���b��N��ȐY��AX�=�ǩaل�B�Oi��"�3RGk�e�	L}>?cp���1���ElM]\�['����q���v��WX/��� �N����X��������M�QF�ŉ���o�L���M���;z�%|Po` 5b
����l;��VX3��նbI�C8,����R��C����g��uc�-��y����0�߷Ё8a�B��1]J3�{]D
����C������X��ځ5�g�%�x濶S
��YG[����;�T
�����=���ae����
���}��l-Ig���C4�2�����<��I ��uQ�j����Qq��,���3 �]��@�Ak'��g,Ç�7rZZ繙������Š���Z��4�����0��ꝁ�p��<S�Q����}?T�9c��oW�W�mz�X���ߥ��t2�/�D��H畍�Ћc
_*��nB���eF���N��W-%j�N~�%�=��?�;�K<��Y�l�?\T�M622o��u���n>�����(Bp�[��J�ㆱ�a�Ar9?XOq��c �t1	sWj�@�s ��IQ������q��d�;ٌ������3@Eƅ��.PG�\�ڶ�����ۍs6O�f��!��hY�%���v��3����d/$�~���Bi�m���F'(9>�\�����R�����--'��:,f�Ҁ�Ҹ}*���v��P������ɢ�΄�b��?���3�/��0"��3u<)��sz|�
��n�r���L�~�>�+�A�I$-+?{�X&�	E!T��h:��6�R�\�^�#��l�����c�z����&�����c����!�;�	ajZ�6{*�O���2É�Y�ջ�+��� #���sB��Ѩ�G�6βl�'�>� q��ƹ~I�����nWR�w'a���}�Ø�����/���;�<��9���s�ъ�߹�#1s%��t�P""����]Kᢤ����q_)4xz;C���%A�z�+%���Fa�N<�ػ����kǗ9�)̂ ��DYQ��k����|&����� ��ܯ���}�F1���*,��v����ti��F�I�sM�[E8���q�ᤠQ��
�w���I�eP��� ��g`ϴK7���L��T��,C)u����l&�sA�uͽ��<�� ����;ҡ1�4�X�PV�яK�'��8y|{Q�*�Y���o���ג�M�2�/
�߹��7�C���l�W,#*y�����L0[[!�q$��c0��$K��.̗�k�IT�w�/���Rm��A�y+�C�J�S[�ŗǅ�X���ԋI�w[����Ӈ�b�OC����z;dX"�?�"��G��Qݢ�0�N�5Q@.�����UA�óv9���(iPep�Su����"�M1�}�W� U��#����O���ؽ��������*�n�V��3�e�"��zc�1�V���	��UF����ox�`�/�j� 5iS�*�04$���lbj
�<L�cK#�JEs�c{vc2S�hՏfU�q�h��}�T�&������
��S���w��ձ�1��_do�d�>T���U��#��<0]�������ť:���*�nG߽n�ۏ���ݥ���7D0��[��� �"u#�Ƃ���Zk?<8[�X[�u�1���s���2�rS��wK}' ��ވ��K7�Υ�B/�� vC�3��n?U�����04??r�z�ӻ�D���w��d�}������u�B����ܯ-��+ף�M���/��{>�ξ�C�]f�7�����bQf�?)���6�Ҝ!��@���]�K��s�Õ�;�,>�~�����5>@�޹�޵
�G�VNo$�=��kx�ӟLV㎹��l�aem�u2�H��Z�Ys�@g���w9X�M�,�j�ʫ�w�8����$�_0\]]�i�*��ʆ�!ЊX���Ψ�������>M�3�*�^���<�P�G�|�B���;5�v��	��׋�1�k*=-V��:oÒ�ި����<N'Sf��'�B��Q�6b�p�<gi��)�Ē*��v�ʌ��Y8]���=
��x*Y 0�663㰬�ijJ�:����n�W#m+����_ѼOh��A³�S����O'�0�~Mӓ�
��}sb�'r�_9P�:|��{%ݰ!�����\A��c �smmN�n���C��ѧdzHz`�*B�9�W`�ea9cwk�H=̉U�HfY�4L����iGr��y2�ڒ"��w��;�_��´�	rS�����%l(�����!�l�3�]ÑU\��=���6�H�D���xZ��E�t�'�m��'�Q1ؖI,� �	�}������8��������h\\\�ҁ8���%�R� _�u:ឺ�Tʆ 5�����æ޵��Z+.Y�Kv�+�i=�$%-���IG;˶�}39w�
��s6&vv�jjj�H�ĩ����¶�$fg ��;*��P'lm��֔�52�#M��	C�5:��|�-�x^���}���:A*�<���.�cU-ȫ�Ԕ$�n�4����o��()�'V���`-PP�_6�|}�+�X�<x��[Һ���)jIyj�|�������p���#nhx�W��mI�蘸d�iF. ���!��N}𢈻i��� ���u��pRށ�W�7ͬ� hO�/G��d< �g�n��ŗhI��jP�b?:1q ,a�I��ܮ�b�$�DV�1����{s�9����*�k��+���2/o�Y�"�$��Ůs-O��3ax���%y�=x�����ϽZ��*?S�+ا�q��@ca��p_���1��9����$����2��7qq�^бd#H`����L�K�C;�W��u��|=��n\�4���:�4�>����>�72U ��pD�dS6EZBl^Q�h�����2��zڀ �E0jH�;#����+�,78D�p2��'�m�]�^{����9�ݭ���( p���re03i[)���[8�_���3d�E�R<�Hc��O.��WV�96Ys<��~��6K�|J�Ҿ��/'����j"��#�w�q0���g)�F�I�0�FGxG��	壙@Z����VZ�DO)�U�,aR�aD~m���[�{���K��rm t�����Z��ć7����?|:8P)ѥzf����KUm=Y��I�}��{�M�Ζ���H�1�J3�FmW�ka�9�k�
����8�>���T�&�J��ͼ�����]ϟ^��5 ?�b�,V���Y��Z�o�o0k��g��O:�S��'늋��o�����ơq�|5me5\u�ͳR�������t��>��7�iu���;�B/����� ��Ԧ��iԯ�	��G��2;�.���J����g�V���&�;��������(ֶS��.�RZ��]�+�ډ��o�z$�M�_ƽ�޸J�c��MHі��q�◺ι�����i.��9'�Qy���6����Z=�{��6%�I�y�m����H�^��7�����P��F��J�~h�B01���l�|�3�u����]y�) /7Р1�J9_6k�<�,$�Q��RQ�"S�F�n�O�DD�©�)��m/��~�T��(��ˑVgh�#��{�� ���D�ǚ���nE�'tQ	)m̃��9_f[ �ƛ��?������slc��j3����*}��6�lF��a�lG=��6J.��3TT����D��[��rҘ����lkn�i�n[Xg�L�<���*���>H^�V�=�9��kd7��{�6�?�Z�Q����lb�^����sDWPl�{<Zӝ�)���HvK;!`y��� ��!�ڱHg_"t�y�}c�b�#���E!�-�b�G��V+p�L�ȣZ<�$&a9������<g�"��;`��7cg�ϭ���B�ς�b�@�����	_T���!N�R��@U�&cJ��fz��\�-��W�˂Ӻ�sD���TTY8>��S'�I�j$�6ꡩ���:���c�\�Uը7CwG�s+(ȭ���\@��ݬ8f���� �^\��ۼ�$�s	�,�ա1A�w��Ձ*�4�.%��Β�5_C4��O������T7���ٚ�,�w�?�@����r�Z��j�������]k��"v<8�I�<��:5j���mO�h��M�E꓌9U��R��tSxzL��f�VV0���
�: %%%�T�"ˣmC��˝/�o�����4�����LD��h�2_�U����u礎Te��'ԷUs���$K ɪ�j�,xy�$��6��[�F�d��w�'�I�M$����@��޳�F�
1�?3��~ �Q�L:x\*���p�aj�B<�����?E�q��wE��K�@~	�6o?�贡�~t����M!�/����V���W�b��+a�o������������?��X���~���Ì��z��)5���L���7�v�kӒo�$@���s�Lx�견.l����|�
���~����1��!�}���6��ҏ;1�oj��C
)z�>E�i�tA�lU)�B*�l8#�gı,����/��
�$Y(j1�5JH��>��o��pJ:�J���`Z�QГ���9$=�\��V!/��ήl�P30O�4Z�2G3<�w��N�ٰ#ƒ�7z+}�l�V�Q�s��d��Q��X��YW1��8�5S�����I��Xx>��M��j�_������_�i���w����}�M�u�c���b9E�"]���j�GH��'Y��ϚGe�PT�Zڔ5��x~�#����1w��x1�c.�N\@�Ģ�Z;v��tA��"���̱	���_����ū����_�"/��oﺘ���V��L ��(����Z�yVN��PN�����	��7o2�,gӔR՗����<i�KɩO��3b�C�kgg��҈a(S���9E?�����3�8D����!_���� �������pU�?Va^QxQ�ԡ�Q�;����Z|�A��Ȭuj�2(�_S�f$�E��w:΃a�vڨ�2p�G--d$��c���	�4�M6kڙ�����k�=��b�9�CB����|��e�n�R���Ga^��W�)��k/�&�9
�O4�b�K�{><���p��؟��r|�F���ѢؒR��n��̂�x �N�	�'�D��6�|�t��45m�;�3k��"<�	��5�����'���#���f�ܯ��\پ�Yd��t���ѳl�*�X�*�3��F�t��L�d;�!W�J���>���t�N�NuR�]��|,I��ՙu@��mx���%yB�	/5;�Vr�*��5
ǂ�g~GSg6w�%Pɴ'��RU�V-�u&�U��-�����4�U3B^����%���Ƨ���IQ.����'U��F��a�,^���)}�f�Hs`o*`,B���	�>s~^�XE2��������=A8�[O%��h��^@�ؓN�[*ZpM��`���)��Cf��I���p^�C-�\�Tr�͕�W�*oؓd�t��"�:�����](�')χ�'ǓqQ�S�G�ߑH�Q��E!�5��=�,��G�X���]8�D�us�~HH>V3n:6�k�!�� �f�-�5�6�u\⾻���Jc9�Af��������	!��]S�!�㦦�������{h1T�:yA�u���o,�}iL�XlQ �0��ӲM�=Ti�,1���8��w�!	�s��>�.�'��|[��ʳF&
"�/�L��9̯�,��dȬ���Xt��5�R��{_~�r�5�%"����*a�B/R8Ē+b�F��9ȉ�ϐ92�Ol�D��k!|��	�_�s��}�5EnH���xdz�����1�W�L�-�	����9׻؉*E��H�x]�n |��l��VN���R��`��_��i��/��&������^d������<����M}�������>HF�0��5����0'�)�]�5]�.��[Y���{�TVM���!p3k��?q�'��������wt(a{63
�ٶ�3g�bX�ߛ���]�����C��� *���R6>���ӡ`�$R�M�@�K0��RB	�mN��XDR�4���CoUtB�V��L�!Eo\���3⬹;�t�:�Ҫ��B�j��k?���E3��^썾�A��^}��S�#�*c���|��W����H��@�I�4�rT�"����\�&:�d�F��&䛴v�{��#O���Xe3%Ҹ�Ñ�fZ���B9GF���a�o����(-j%�IeeZ
}��v��n#+�#�j��Ӗ��gL�U�>�4�8��0���7
��DN}���Ki>������a�zU��:�B#��-�Cx���V�J�6��P%�Y��5^�R^,�E,�_���8�uS=���`%G��ͯ���~I�HlP 9}e1�;��ڬ�r���֍(�}��L��K�u]���TQ��m[����G_��9ș�k9~���y^R蜡y[Ԙyb�6H�v��2*W���Z���X(:|
ل�������ͳ>|4�U�B�@��S��n��@��G�iӟ�� �Y�J�3z*wx9���x��X���e��>�ұϜ�8�R �`2F_���5G�t����R�\@(�r�p����@|�?^��ksO�"��_�W�ȳzo+[�nב����� ��OO�@��Z�p�6`t�����`��X9����d�!�	S�'@�y򭖖�U�=�@���%Y�{a�s��|%4���)긆X��(QÔ-�+����8f�CG��Et�k��=��1&|��ʜI+���ߞ�nn��Y:X~���|��b2�.rGk����.��42��ï�OM�'_��44��5��m1�oc�.�+�����6��D��[�R�q�Ѻ����y�S�����..@���Fp>� �'#�]Iz��k|�f�����>�wf���lc�r�_�h#���V4�J%�/j���w�ף~s9 ���DFps=�(�T�P���A��f�V��S�6-�KHap�$&&���#��۾~�+K&��T/K�]I7n�� �8�WQ�0�ǔ��qj�5��X���͒k_���^�QvKJ��j�J�ΎL�6�����m�����S�[��s��]b�%Y�=�٢]�UT	���י©k��):����Z71GT���0���<�37�g�Me؜1���jv�s&�ͯ�2����y�Ȗ8o���%��t�9�~�j�#��G0�����Ƙ�P���Nt�\4�BM��7F_a��;���N����jܯ��}\�e��YAR��t���f����8���G��C�����M�0=�X����Ď�W��J�k�Pl{F*��bxK@��աz=5�c)��Ă]m�ֹ����<��""�ߋn�z���^���²'��������m�J#�*����$��:��b�Es��74�LH�Q,[љ����	����
>OJ��p�0EҶ�9)i����	p�?��2��J|�k�;z��*�?��ԯ��|���& V��ߌi*�\��أWNV�@�����[B��P����D�"�����cE�B>h,d�j���}hO�R�i7/���٬  ��b�c���"�x՘F�/Yp�&׽�q}���]@S��	����{B��T��h���;�Y�� ��)�Rb4��٣�">۩;�:�h��ַ*�^�]$Ӧ𾆕��y�|tw0!9w����������s��4�r�Tg �)�o���m�cHs���g�F]2��P30�j���}������b>��y�i�g�F�|�Vm*���	�趝&�R�XEXqX88���A���ʹ�*j@+�
!�j��g��DZDƯ���D�W�奴��ݣ�����ԉ} ���}(�s�S�O]Se��}��TN*�0U����W�4�_7�|�o!����5&�����f<i]�,�����ZX�V�a*7n�~P �|�]�6n#�Ɗf�!���@�G\^>���g�b�'���2����k�On�)({��gyFl�[�"X��SPRԪ�U�I���ߨ�,�Tkܚ�c���QV$o�x@�m`� ϸ��U��4a}��/r�������Xf#��γ�'z�$���V�w�Q�i)S�O��9j�0��O�=h��!����82g�+��tB���>��WR�����%9�{EO,sZo�S��=���W����2&[�!D<<����f|�4�"�B2p3z�v*��յ����	D#��H*�p��E�6�Ȇ�꤁�i��#�{�w��x^D����L\���Wjm��q7�+'�)4Q,��o+�Ӏ�z}	i�v�G$�v-�%��o�;��g�q����:�f��Bw�V�r�?���#Uj7W���)�K�A{��Uob��eR/l!�(���\c��S���ׅ��L-FYF��}�!2?�Pr_\���?�[吢Z��fަ��E�G�iw�F�YJ�ɚ	(1���8=�����oOC�T�3~�[63��a��j�Y@>����ym�EA+a�������H��oiFr[~gL��3�/ya�lŎ�����$n�?m��J+ج���qS��~�/i��$g4jR�Qد����V9����pm�~�P!�C�38Z/-��ejR��_Nu&�����]�7Ga�VQr�v���81&M���[��}T$bt�G�y��=y�����˲B�����kv��H��]Ӟ��2�,XQ���o�APb�����ʴ�~�Q�{ށNl`�+\;*�!f\1�38���]K#u�Թ^xBc��\�}����
'�*���#1qv89�`+��
Ao��)����X9�������v�!#���)�Nl}4�Q&��m�&�X���0`1	D1�����})�{\���~�v�B��(�l$�1R�DUşQĪM��F!*�jK/�5���� �p�+\�Ny�۟	�,E�j��~0|�t����]�I9�Q������mv��@�;Q	�_�����>�1=݉�x&��.��|���M%��TJ�2
 f|ָU�6>-�4:�'c�(]�I��_����!O�zq\.����pz�3b��z�Iv|�O�!0S�[�';��"�
aF?o��V�m�T<�F��Τ����y�h��%ƈA;�͖�jS���^cf��e�&̋(5r�����l�Z����pk�⾧d\�ˌSa����%A5���>W{Ed����&��:�U~-�]�xBg�xp��V����Q�o�1&.� #Q�GΎ�q���w�c���w�$����ܮ2���R��Rh�h"�f<VZaO��c��uR�ᷓ�9�	�R��J�7�Q#]�+hU�Jz&ֈ1��&CQ@v�]h���T� �m�Jú�p��>�:[i����c�S�`~ٯ��#� �`�ߐW��y����Fb|XRg�w5'�bq5ds��3�D�s�@�͋�s���:� f�p �grd�P�o�9��B����M��+r�z�D���!a���s�>��|QK�L�%����5�+�ب
�cۺ�Գ�
�ݸ�FbY��NI$������5TH>z]��=Z3���4���o��&c�A~�>;l44�vQ��z\�w�9$p"垯�GM2�Zb�u��־.�����H��F�#[�y�L=�+�0�`p}� 0ߛ0d��Ŧ-�GlI*`�x�M�7l��/= ƍ&`�/��'����'u@��^yU��`m)�/~��ꢎ��p���5����z�XA�]�R�T:�K��g֟������j\SP5�#��V�Ҩ��uR��͘�zV��R����% �B�E�k��>����ZGSL��WKIk�3�-
c���������#}l9�o�|���Җ�'��s b�]N�FC�,���Q�-�U��y)�e���\�u�W�l�f�ږ���zOXK�������A�#��ب������Tt�@����f���ȂA2:�f����gD�5����#��"j�,j� 2.��7'Ф�7Ô�?G�(�tCi-����B/�5c���tm�h��Е4M�0�g��xӗq៼��`��p�$&QƊ�*���$��eԐv��y���Q\�y��o�� �"S���Y�vf��k�R��`67�c����?�����9��g�6���wR��m�̈�0�&?��*�TP`�ǽup5��+3�"+�t�h%&e��/�@U�+��Zc|�:üz�����O��NF�y1�[�
���-�xN6��q��"{���WX��nb>�~|�Sw�P$E��p"��(%B��ME�%�馭�37C[�ʪe��T��\�,D4���d���_0${��������1֦"��Tћ���,v��\T���1�E,	��ť1�vhԉ�'�>�ۧQ�h��2y����O`�����4ՓA08\>�D�l1EYĘ�nC�_i���	?��s�9:�`����'9���ҹ��]،�_tb���h��h�r�cY����+���W��X�C9M8`����u���n�����m)J�N�I��FCtZ�O&��l���ϩ��,�^7tሴ�^�ff�.����cw�}F5�1#����Ɣ�L�O�Ȁ�M!0�3!�:I0QHy8^����M�FE�d���7x����7Fn��a�}j�?>a����F�Ӎ�wχ�+����~��o3_�9��oh`ȡ��=:~+g� KǑ�E`�:m%>�0�;4����;�(�|l��)���3	���~;�v�u}���q�զ�EցB�UO�ؒ���z����{JLJ0���%Lʠ��Y��;_���gN}����uΗ�\��]�ɕ�~�d��㛽Xi�AT�$}�7��Rҗ5�� ����e�>ãm%�m�\[b��r�p�[鷻B��7N;�<��,>��;�>�����M��q$dgo���8�
�X�m2�^.ĉj;i��w_f2���������R���2P颥ҮT�����ڼ<����P��{���ę�le��v1�j���6�1�!����x֘d���4�ܦ3J�F5ĺL�]4d�z����n�
G��Y�'[��$��R)���dB�C���2+0�=��	ays�ygXu�x���<_l�Q�j�[���u �x͙F�9w��7�ϡ�5�����p.��rl7|猽�`�� 8F�����'b_c���U��F����3�dd����y�{;���益?��SJ;���-�X,�R��K5Q�������@�����[*�epe���%�9�[��L���Q�tvc=:6frvC<�������0>�˶�`x�2���1���`�6{ �+Vع���r矽�����7�j]wʜ/�J��������_:b�N�/�˶�L8�Ie���a�K�<N�0 0�Tx��İ����H�80�W���L�u�$F9��r�	�}7��r�/�����~�w0��\�%�f����]=��<�<���Qٌ9!h)�P(#$�n�p�r���G��@�
��n���<to-,�!^=O6N�R�Y��~/��6�H�	�G{k��g���=.�D
M��7�~���d�V�ηsZ&��=8~[(h����r�/ҧw=	` �X�v�`G; ?�aLv&��1�ߧ��)<|���u�x�:o��
wͮ��-����ߛ�] �� 5�\�
E5	XJ9gt}ًf�W��u:��� ���\���\�ӂ=�DnN�T���m��
6�Z�����D��:�����I��~{�� ���3V��N�A���sOs���͡Z�?~��	D����6|�����ړ�E0Ձr�[�2GT��).��{"�rL3s2����߼֐��r�(�s�G�-�m���V�ާ���?0�6��2J��~�=�� ���9<�1���qٱ��p9J"�9�ݜ&�!d�C�J����"`	�}��E

ǡ��Δ)*�������X��^�ʉ����_i���Q�ݨ��l��1�3鸍���[�MǍE���i"�d�
�|?�0YrD��@ր.w{R�d%6Z}�`m_(�1!��԰I�����,x�M�X�ٯ֡Z�w�k��8f<ýE1�fr�i-�/��e	l��Ђ�_��h����),_v��y
�H��b�vt�[���j��e�y�M�n��F\<�m!�eM�cD���claY���าv���'$'���H��'L��tWc	�$��N�)����ai�B�e��#�[�O������ԋ�|���3;dly ���{�%/TSe�QV�C��T��������H$���{�/'.�L���ar\<�ɹ
\����V�e���0��cnT-5�s�dR��h/p�Ӭ;�����'��H����gFD������8A���|j&�&4'0�&!��DW��%�a��u�}Y�6�����T�c"0Ys��z�<2J�
��Rm	�����B��L ��/��9h�����L���Ϳ��������/DtK�.��{!r�9_ZX����#������a{v��I�|� bϦ��E���p����4��#�A���ڗ��1i���SSP"�6,a�HI�#�ϼ�v���0�pM�T=�HXl׉;���ʚ?۝�����R"۰( }!�G�F�m�ٿ�-$���_o�;W+H�CX9��nm��2u�"�7��bu�&󞏥f�ಪ�ߑ@�H�6m�T�Σ��.)�=Qu��($[l���B�,�?�~�9� qk��VT;�A���?����Fg��c�͢螓���ǂ��:�(�.����W�7҆��9�����w����������?%��&�Z4���t	��E���?�bB!�����q��)l>��9	V<D���׾KL�&Gm�y!���o��h�	�JcG���~�o��E�s�
��:��\�p%���/��>����-L�h��é�D�w�UM_;�c��[���Zs�GA��:�	��R�S���������:;�?>��S菤��_jS��U�w%UE�^����N���ooe�Ԕ���h��%n�m�J  t��{,�����5������&a����k7���5j&����R���b#)u���y@q"�z~K6�T��b�UE����)JH��WS������Y(QÖZ.G�BS�5|�`SU"�?R�̱�5%��U=J.� V��Cj�$`��Hǉ�c��n��7`.v����(�J������c�"zH:����=>|n����ſ��7C�"u�6
Po�u�\y<���G�f\���ء ��2�O1ݪ����du�|ۘ���;�5:Ed�����h�hI��*v���l�1m��)�&�����N��=����ML=nl@����xR*O�ID�?%�L!����W�e�%U=�-N?�	�4��Lr}zV9��4�s�E0��b���!��G�V����;F��v��D������o'&-��)N�v�?A����6��D���aF��%U�<�m��� ����t�N�F�0�e���s=x0>d���x2$���� �#�@�7
ӱW����3�;�5�t�e�zD���ˢu
�˛��ǵ���38K`�W�]� �_3��S>l>����T��$lo�ö��i�Ou�-N��__��V��c�љ#S�����P�����&��a(q)m����K�gH]'$�)Ѻ�h�j�����28�*��Ҹ$�	Br6��g��8��?��������}�������O?���A�/��'lˇ���B`OD�@l���O]�d�
�(17����ed�~�X��&�$���0	���-Fk#�G�]4im� ��l�;*�&��� X۾��^c��u4w�S��x�CU�A�!Ǚ``3ciy���I@��A�3�#���鮈0�a$8�/��g7$�[8���A;��#w�?>� îpp���Sl��sm���s�����vCZb����Qr�d���T?�TA-�L%� ��}�&��9_j���>t�s�OQ��,��P�`zS]�$lZR�4��*�0�,o���C%�Y�jp�	6�}���
x*��=��s�n!6��h!S0��U�4~n���xv��{�e��k.^��+|�L��ׄ����9��y����YQ�稜�]G��.�
d�e}�p�O���T�}gyku|"����D�$\�i�*��g��(�"#���݀�cd�.��G$����F��l��ęPO�5zRk�G-O�I������&����lXH���$!��sǙ_���8���%�u֋�x�Q���_�d���u$�{���:�H�����ʞgȡ��V=�o7k���BAT��	BI�e�;���d�r���P4�L5{N����M������h�yA#�ֲX�,O�-I��-�m��~A�2ml	@��RK˰@��1Z������J��� 3b�H��ն�RU��k��>�e�W1["��6�����>Z�?FJ�Q	�P�@�g��z=>;չ�u�L+q�f�Fm=�93씌Hd��������a�	�+�똚����� �ï��6�P:æ��D�c��{PP��'����&��<��h�P��,$0�Ս�����m_�E���+�����n���/k�y���62��{Ԯ8);�����<�]! ��N塠�В�������ovY�����ч�r D{��ɋ�bX�<{�"m"�'B�%:�Q����y}KY��.=�[L��U��V���M�6�43��u&*��w4�vRTT<�	�}JM��2�/fff��%��t�.�|%�7sV�q�q�_�2����Q�x���`ᛝAOI�d�p��0hn]��5�H{eh�5�7��b�Sޡ �}�˰p����Q(�,D[}/	�;��.b���O}&5[�c����zp�y;�}l1��u�'(f�1;r��k�nGϪ!�;��^n w���d��;�S���׺$\! ����C�����&�G������]�^�)���ǘW��J@��]F!��_����4����M?����7`KC�-�$uY2���~Փ	ȫN�x�3��"m	�ߡj=�mOx;��%���j
�-��)k�(��]
X����l��t�ٞfo�[��9�Mdd�3�!���/J�`�B�l��L$��nVy��[��+;&+�Il�%���j���*�%1͹�	o�:���ۧ�ڇ�q��DG	��Z�q���f��.�:5�}����F�p���w�J($�)�,=#��:���Pwh������2�`H�m_�&xk}�TГ��G6���2�,�c��х+&ϻ� ]ˇ����p�.��$$���g�^���n�����a�ڹ�sx=Ly 鋵�J���GM�ɼ�2������{8X"
8jad�*z3�>J�jR|�T�ھ�u�;��pE����Rel�:����ɏ�Z�������Q�%8,�b�T{�dھ�9
���H��M�+����{��������S�.=��>���Li�ΈlFň8-M�;���NgN�g����,�s��n$x�#�4-���\r��Z�#:>�9LH�C�2�r���^��a;;�4��g��(��%.���%q���M�oL��RY��T�R�ui��ƻ��~˳ɚ��i��n�m��Ծ��25$ȏ�/T�J����W�����j� ��Pw=�l�T-��l*<�=ʰu�^-�-N�a��"�u;C<�����:�J���c��H�5�	�(b�R:��!G�zV?N��џ��w��+�'Ͼyz��߬p��6pR��M/(UH̴�/_��;�<j>|)f{�J����O#)�����\�r܀�,�趴�t�.�G	�߽��\�hSԊF?aaɭI�$#n�#zC%_�*����Y�_
�����7(�,C�U���C�>�Yʯ��o�'���f�N$������Y�S�̱4|�����K�E-8���9�m��ف6F��&#�o��>���Gm�c�5e�Vn2Q�����^u7t���3��U��4<���b�@º�ȑ��ai��l��%d�N=�\x��UT�)��`��s�zX��ʍ��j���[<nha��j�JY%�_-<ܸ�Y�h	�gn�{~�F��w�Z�+$���BE�¤CZ��E�8�9gB�`��R��#A�l��k}(��_�'�<3����������� PK   �	DX���7z  �  /   images/be8de2bb-09ef-440a-a2d8-19619bf9d0dd.pnge�uP����iv	Y:X%D$���e���T�[@���f)Ii�R)ARZ:�����>����s�g�{��3��+Z]U���PA���֨=�A��U83�t�7�@C���o�����B=������r����p�A����|���ae�j���n�u(J��FK� ����>�&j� ��"�>ݽ���vЦ;������p%̑���a�Է���Z��R�P�Źy����S�3�g��'iĞ�j�8�Z�%�Ww�G~ڝ�ջ��\1��pY�ӭ�Ǜ����L�>�����֣�I�'99y���������_�_�"�m�g[#�w�G��,���o\��%�*��&����o�i�7L/�f��;��`�Ҳ���>r�92��{�H$�s�٣���<??����QИ���?��)�G��5���>����7��II8 �_��ia���0-��;���>������r9�ﵗ� v��eE�|R���k?�-?=�l�o<�Cj�A��Ӳ	~�e�t��w�´������K(�
�\���.?a�D	�:����'@7ݬ���� ߽�����}aG��o�d5�J0�#�I�� GD��i��p!�X�x�l��G��@j>lF{�����O���`�'1�		��`kQ��k�n�+�߲֕VR���@H&����ѩ�_Ĵ��� w����[Tx���F�s*�m�E����N�*�]cX|�<���"�P\��҂G����ؕO�i
�=I�Ҩ�8��#J�h�6:N/-��ڇ�-N� 	o��Y� �����O�E��{�
�/���L�kp@�wy	d�Dލ�V�����M�O�ru�Ñ���7�M*�P&�i�$g�P����ơMؒ�?J�x�]�'6J-M��%	т���bq��6K*e'竏*��ӰM�%����[��w2��S��፮E�@y7�J`:��;��Є�>�L�Jq��1x��J�
�O��[y�mN�P���].�H�ԋ���k7�ܢF�G�u��`�e�Q����<$��v��a]A>4�6t��J�`���&���7k���sJ�=%Nm��	�烥��+g����\e�tC}ە�nsߗ�բxy9�WW+�IfQ����ȳ�ID����)t-�=	�(Ke�z��+O/L8��0LDQ6�P6�(�T8��C`�)��ڔ|Ox���˧!Y��u��`���8���[�}��f�/�\��S���8�\�����^���B���İ���B7[�2k�L�t/Ũg_1��ǃ����p�ҌI[�A\����&I��ϸ�G�������4�ihI�	CX8`�<!�����3���xnՎ}m�}��Hui�!�6��ޟ�^��D)��_�]��� ɴJ�+Ţ�ۅiiC��
_�$���b���BF�GHā3�%���㘂>�{:���,?�f=�i���$Ga��m�Lx B��Ha���8���݇�ǣ�4_�(U�&���fY-2F�'"�A�^Ui鱋�lB�!具�"ZX)��חI���r�6�9y�@�nj��Y�L��KvQ���� 0c�'�[����ǘ��1�ߔXb� �ٙ'�x�˓�q�
�b�������Hά0�A�8�.���nc,��|qrZ�ޖ�����+Gٽ$]�6&]��L�u/,d7P�����O��4��rtQ(�U7���[PX���Қ����t�����cp3�
͵\Q���l�;�n"�;����p��y��!�;����Zt�f��>jg��ƾ=��O/�^���TY�� `#o���t�L���QD�����-��}��B�M��es���wh�Ϻʩh3im_�6Yb���lc�y����]�0�Cw���0"�M�2n;��85{���Mݱ7��uҵ`|%A�z!}���
i�VT"�X��e>'�}�	ռӲ�H±���l���b}�?W��qɄ�������E�W�M |��L"�!�2WW������tcPh���wDpo�F�P6nh�����[���a}��I#{^��X�p��ŌN[��j��*Q�==�%<2���;,r��$���7��_�k��ƚР��
ݪ�Fs�S�}[�|W�eG��������~�n�"Do6�K��u%����a�E8��F�D|��2��C���5�^��q������<O���ƹA��s��(��4��(gp���9U�0���޳���TTFHQZj���z�`�k����	Y^�-e%�ˠ���܀Û�����Dq{y#�r��G9�2I��"�Ke@;WҪB�y���hF�z��TL7�&�ȨD5�2K�> �Z
8�OfQyw�'�!�2�q��-o=lq�E�O+�˭�X��'n{�^YOI���v����y_�V��o��)�\q3?Kf���^��T��l��]�Tӯ5�Z˗~q4��#���W�`�����Z�������ed8>%�Y)-�	� ���'�;���$g���)0�Fǔ;`K���l (���y���S��O��߼�>��r�sQ��l6<njڛt�!
��<[mg���s Bude��g����1�\��"�}�&��2?���'K'"��/$b��o�2v��j��{���y�0j��C��3ngZ�;�6�`�ݜ$;��TJ1>�jll���8�6a,|��F�]�ٹ���۟�;��V�Vqנ/���õynG�jo�M�+�ݧ§��~��'��I�4�^O�����H��/Qδ�!����jz3�����͙�b=6$���nE�{��k'v��s���)���`�E���i�g2#�C�=Jj�MO2�����z�֡�?h��F��8��y�&l~�R\-h3U/�q�������������K�h��|�����X�I��r2F�54H'��O#(�Tf��*?�و�����}��"%�����ۯr]�C{����T3����0��6��{�Z�h=��~cdr�go��Įj����g���3���f�z�g�[&�GՉQ[. �WNn�wU�o.�#P����$t���!� {z�ѐ��s��L&�_pgk��d3��[��]p��d�*q'����wUN#(U������~o�0�����g���J8�rC�@g��%֤K}a�( �؍�Vy��%V���(d�ru޻�����q;��]�J�W�a�~�&��L3r�a׫n(*��l"9����t'0�@�fE������t>���Uen7���i�3-�7Hw�Ol��;�����L&L*�qLoFJ��?dǰ����H[5^(����+1$=�\���e�9�L�^�^b.s"vY2�j�|�Z��6y�n�J�E��j�i"�����kd�|��"�a� ���J�����B�F���4d뢦@;�7T�K���a��x�Ǆl��!y
6���	�,QjK�f�3�	~�X�)X����K�[�h掲�4O Ϸ���V]KV2���<�/�pn� ^N���. )��r�׀AᏉ�<�C\Á�}���Z���G��ˀ޺����v�N�"�W�ȅ�؊���ʎp�&{������*p��BZ�!(���������(�[�S�13�i��"P�%$w�Dd2c��[�k�Dώ�ǚ���ux������`�����͇����Q��
�4�T�f�k-���;��)����^��Mc�*���ggҊ�գ�n� SE6N��n~�iP�/�[q���ʮ-v܅y�R�ˮ���뷖�����efx��C�N���ɽM�O�gq.?���ֱ`�ь�ăz��'bSrԍ����to�7#���F�a/�C`�e��V����^ZF
]~p���6q��$r�`��$`�@��N���y��%5���#�P����ڬ^�C�q� 0��)S��2p5=�����d2���g�Wb�>C�&���]�Fހ~�Hl�G�����!~�UU�F4��魕��]��#�rNWN��r�~E�Ԁ���x����ݛ�:SUB�+�*Al:��}���P\����1���C�uRO\�K��X�}����6�be�~�ܶ�_�x��8y�iL�L�\�^�܎B1s�,<o'��=��$<����(�a�8[�B�Qe��c�3��4Y�Ҧ/�u��	T<?�N��F���r��|~��6X5A�H�;��5mЄ�Y�޴�m�A�eU�9���VtU���G��{ؼmX��6���tT��J�m����e�x�4�Mۇ},�n2�H�.E�����ʥ��Ftv?���f�[��H��.Z�;9j�Z�����t��~����e��V�K�*ߎAq�D��,�1TP�Fm��c�
��z-��]����6�eX�������l{�U�=N�u\:�M���]M]�T6�c���(��:<&���!�w<�q�� �F�s
�6� �`��|ѐ�
�����L�����qbЏ��1w��;�i ��7:Ќ�_�?����B�{���F-�`d1AcQ�o,�b��Y 5�d�{��A�l�������;��_�U		'��=;f��?�U�	��5�|��������oWtp�F����t' Yi���g��4�L\C�[�r$�	n��4�F��μ4�;h��ޫS��W[4�[��u�jX�>uW����G��ٯ&���ۚҗ�X9�?�Ur�<�6�O��'�[�F��_^Vj�)7c�1�z�s��0�����oRrNq��t���f�8_Q��2H��q$?��AY�j9��p�_�{�U�6����-��DMn�u�z&?�ϸӮ�dk`��Ķ9��_Ā��iA�5��yv����ꋶ���M娖~,.��^�gį?����J�a���%Yz��v��#K˸�������*C���}�Hx�ټr:/����\��,^�A�y��n��k����>^7�t�L��'�
D':�ϒ����/oٺN7�]����}�j,)Ѿ�R��ɲ�<�2"���	Ym=�pXG��-IgN����KT�lukL�>����L=�Z�zAC�D�F��VZ�q*��'��������Zd���6��7��g�M:�7^X��Z���h�!��Ŭ메"X������x�9A�6�	��O��4
e3���h��zDxg?)��Y_�(D���,49�jN$��˚ůE�C�	g�Qe��f�{z�0j�Nr�̡�9�s?j@Ǳ��Ml�����C\�n��{��9�ۡBھ� 
��t}����|��Bl�t$�#7��57���~����Q� Ll�d��ͽ8#� �1S�_?�1p���������-�JZ���]N1�Wߗ��9�pP���@�?Z����3�U������H]�'��(5�F�kx�<�@���qbM�qZ���(�����|������i�A�n�<&D�V��̒���x%0��=���u���y���h�����kӶ���K��v����yMc�t��8ZvR���֪z�~ń'��rb^����w��{�$� }�i�R��*|eciN��<`��Z-����0�U_��e�3���K�s�֠W�]�M�%�hh��)����fO�3M1��b)��?�]��l''�M����sTBKӨ�4�׵�j��
�����9y��ऻ�����j~�iF�T�M���k��>�����3Wo�`A:�FH����X��p�>��
�/�ii̮����g�DU<�&&͚��L������,(=��+F�:�E�,�0]޾8֗+�_<b�|}���u����X�^j���cL��5�Qb������Yytl��k�ǨLM=��?�/wĉIX=#t��qxG"t#��*ΟY�]�t��7�1��_#җl�U�S��q����d��g&t�znn\��{,!�)B��q�P�P��p��K��M�	��޶��C��μ{B�ZHR���x�X�OS^T������9�x�sS��$����R��ǹB̬��F�1>z|65l����M��h7,��>�ٱ��2�۴QBb�(9Rz����ϲ��>���e�������%�z�8(s�IS&�/hDu5��o��r�%(Z�
���;�ρ@�S]��,R������ڬJ��@!�_��4ƒch���%ѓ^R�6ihJV��٨��{��`��t�\FΥ�E_��+�le��_�o�E'��V�MmE���B��������5FClwh���&�3�;J�K��X���HM|ląv��K��D4y��-��������[�V�~���<Ź�@����7�:I�j����H*N�W%J9�P��O}Q�Kj?�Ո6l���>݉�g�����r	^�S;�~;"���Տ��z�n�f�2�����XBDF�ڦ&Fީ�����>{��58�QkH�';�:�1-Clx��t��i��)W�X
( i�ޙ��2�Ow��9?�׏��0�-G6bdN(�����7�Y�~�{l�vz�������mg5\�#{�����0�N���3������\F��7�H��rTD3S�~s2������:`�8�ER�,�;��[���mtܻ�ݫY�!��w2CS�ܻ!�>vK`���Uf,�&��xH��,9]��c�b�h��R{���8o��K��z���
�y+I�Z.t�Ӽ��:q~W�Pzh�Ֆa�Bɻ���
����+k�]�|Ȫ��H�U���5{O��ǔ|�I�͡��^	��Y+N2W���"�S���V-$�{)O~�����g�;5��d/"@���J��W��txnh�EU���Z��.YL��<G�3�
'��!::�'�J��؉/�Z��F��-1�͸��>�������M0BV��ہ#ׂו!����|���D�Ko�<�EY�4J��mZ�5ԓ�n*��R_�|LMܫ�\�Xr���(�bx� �(��SK��t�2�|�x��]5�Ey�KI�i��c�A���K������������=�	����h�U͡����*�f��� PK   �	DX$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   �	DX$[��>  dy  /   images/d3938c88-0382-4189-a86f-3cd234ee676b.png�XS�/DEG�3��F��"A"�iR�Ch!JPG�hPz@E@B�5DA�I/��ZzhI����y���~�����s���yx �w�w�k�k��Z���i���ñ ���+� �}����J}�n�k��o:� W����烞��} �z������@�j�k�p�E���A�Pg�=\}��z�?��vL�k�@~��\�t�?ya$�E2*��dر:�e��T����wkn���@��Y�G�ö�7͋�'����+��Se�o�9s��T�Z�EFl��G0B�n��q?i��~�m�}{,�Z�ô�J�j���Vf��ʌ�Ǯ�8��|��_߯��?�ҋ������`Sl���-Z��{[U���Oe
.��O��|��5�׉�V��Rr���u�g8b;S�p���a���1rͱR��E2��ď��&(�|�ӡ�.�HQ��:�|�_ߨ���*�7?�qk_*��ʸ��~��r�6�1G��q��qt�:Z�����@y�܏�)��sA�{�G=�x6�e6�`y��y��>�)Wbj�}bZ��~�=;;c�*��X>��@�M��_��#2L�K�W"1&k��c}�DXd�g���yJ���}��U�;����)���7�腳�$�/�Ē�5��`�jn��6�x��0q:���7�#��裦��c���ޯ����y�\�4�q0�x���65�C��Cg�Ő�V(S��!UsJ��!W���qp" i�����j�K�,��9�ρ�MH�|��&��	�`�p���V���O�����ga��[���u������Do�#���x�-O�QVX�bK�U�L�L�9{�5O?,��~uV��]�%�������?h\)�Ȗ�k0�`�H>/��+r��=�*2����{���>�
.��ZX��$/Tn�S��3���|{y�p��������B�{E9������b��6oe�m;�J�C6K�7J�����J�X����{��E�9+���zb���&ƶ�{rڭzSN��&d����S7��c�r�԰���(��)�;���ܧ�'���W�v�
�3�tڐX.�V��E��H���S�y���A�����o�����j��>���R
���U���������Jv�S'[��tB�\r5�io�ȵݲَ�	��-�ha�̐٘A���$v򱎟�&J-$W�6������2M��[�:����\!��(�jhp\7wi�ȭ弹���\J;��@pl���	:Ӝ/��%t��**n��/���<���)��ؐM�y,��#g�Bóz��w��
iB��j����j��:�Г�t$����������p��+�rs���6�j��Ba��l�Sݛ_c6��t>"m�a&0k�\*�Q"�pML��+�bv|�>MU>��B�r9�CG���/z���儐�̽�|��;�:e��5A	�d�N�olC7��bO�?����>b���МQΉsCoK>�,�٫o�ٯ��^����TOG��X���w��O��L)�:t�"�Uq�k{��F��w۪�>0�%Ii���Y+d{<��3S%q~�=�Xl�<�!%��0[K6u �ʯ�;�f�o���ϕ��X���ZE�����\��m8�4�бy��d�
&DQ���F�k5��j?�
d_��#F��l�r?)�Z��=�ya�Q�պ����=�^�xY~�.���N(U��P��p�}0XJu��/�s�wX�QNz�I*�M �
*x��Y��6y$a2P'%ebI�C�(?�ADǣ�� ��eS5䗖��7;���&�?����_Oh/���}(��n��c��:Ir8.��J^�@�m+6�(2{x}�����6i�S�j�sZ���!�6"k�m��ǌ-ϣ8��B!���}]��3s�s�@*�o��4BdM�hx��n��T����)jm}��Y�R������@H7p�X*����l�:�}���w
Ka��+d����,�|`q�t<{��6ܲ�^H��\�����5�,�R���`ڔ�_��u2㈺�{Q�ʱ97]s���o^Ek4�Y2�Z(9eY�!tf�НW9S�p��$���@�ܙ�`���T��l^�w��(Uq��ʥ�ʞrF�# GE���p͝2w�t�������o0��#�,�@Xp��sU+�
"s6�au\_����I�~�5�<Wǟ��8�X���Z���3���,��X��EA�s������k�\�Ќe!ێ��M-��~I�M�(�<��IǊ�UW�嶈�y�j��O��lз�;�6���*�?��� �L�a����ڰ?v��및7������f��:[�gW�X�2	�����θ���Y]��xkRS�����܏@ y�4��cb��ℤ6�h|���6��R�-����a��hǎ?�+�=j��Mַޞo5nz"`Ϲ�*�Hjm�#*�B.M��k��q�uEǃtE��F��Qr�WTƷ p����!����g�Y����{>�y!�7����u���3�P�!U�*� )Vj�t�U��S����[��Cm�]�L�'�_
ǂ��p�h �B�S���T-5�XJ��X|�+�x�`���o���Em�u�w��R;I/�;��kGae�~�/;(l�u�"��ʾ?��Zڷ5�6�b���)Ջg4�ƔDZ��Ԙ:���Mh~{G/.p�����"�WNݩ/��^�M�R��[l����o�1Q�oU�ݩ8��GV(�rƬ�WG�d��MS�t�`�Ԉ{7���vTQ9��]�H�U��s37O�����Va>���K/����BN����Q�!�� ���#�|az-��?�SX]�r/4�Qֲ�����#M룣���L��}��h�[!/?���<�<�T/,��.�hOe�}�ꓒ�Y�p�xXy�3,�7er��!KL���c����#T�̝=�O<�"e!	��(���{ep�_3ј���"4cOJ�V�$J1��!nğXحe����Ap�&�Hh�I��#Y�ԯ7OVN�em~aJ|��Le%ҽ1/�!O��'�NF�	�L�&���&;1h"A��7u�i[�W5��X�<�B��
�\���	��.�p�\�p{���%?���x���xuS5�ɏs��ӹ4܄����+E�)>�"'E�͙!���w&�A�=C���;�f�j�,Nr��h߾F��{�h�D!��8U���A�۠q�w7+��]	����^k�&��\�KG��,�h�� ���1;2.�,�{���s�N�/���@9u,�;F�(x{��Y��Z���;9b��wkG�J9KV F������9k1�����;�5�b�v��էsY���'q��Po���ހH���|��_\�Z�	�[��4U�9NՇҀ�['V��E�D�W�F���z�:&QS��0�cA���,܎�~��Ԧ��!
��� �f߹ia][�����A�M2V���KTA���}��p��h��+����0#|f���x��v�	�KL�"�_��Q�s+�VRl[R$0�wJ�N�f���f7VQ��d6�;��ݐPI: ʍB�uscW�"�	����<^��2H �@��Zx��X(�7��[���X�A���Q�Ԙ��C<�p�� C��5�"T��-1w��Pm
���{o��Or%D������|]N��#��ꍴ3��X�������r������v���8��x�"p�u�m��B���Ҷ8�rm��C�����r�4���}�IGsH��Z�v��y_!���cs���#6>3�ժA�&l��u>-�6���^�(�}�י�KtJ�\I�A�;I���j%`�P����';.8�6G�m�<DN���6�l�Z�pYʍ����c�����b>~_�k�/|��I��1��E�;H\��y2zA2yqd?^���:[��J����ſ�I��.=��I=�~-�\��A��ҵl3��b�r��~�v��D��x�+�5Ǆ�^�3�����;ue�@e+.��N"J��#͹���t�
pS��˞����t�~�d���Z{���~ِ��e����n��=z���}2�aE)��-`�LsZ̅�̷��1O���m�hn�k��;��ivA��;�̴���`R�Rɀ�M��9�����,���[�+���1���2B.r=���?�����$��G!]����a�/�8Zi���[���1r�c�c�xm ��8H�ԽrR>��;s�׮�Ԓ5P9�(H��ߜW���^I�����B�⌯Q�h�5#Wg����J|�����5	�<�~����
�R/�����	�	��^��m��v� N`H&�?�W����=�~���`ҵ׮��8Q>����)J����X^|u,�	����u~y{9/�	���{����,Ч�3����=4�=ي^��_��� �r���3����o�uw���l��C�5�����U��|MP��ݿ#?@�n��O�����]�Ë������-=��5@qq�O\]�-��<��u$ew{���Q�)�V�$�ڲ^~�?�Z�"!���)�����v�."l�z=�e�R;NM%h�1�3��U�b~j��|�q�� �E�@��ȅ���BjX��A�t�]��?0��E	� �b7T�:�dWk�-:���~����/7ȴ]1{�% �$�ɦeS�8��k(v��v���H?[E�@$&��H��t�>1�v��(H�HG�]�����c���wB^��j�-�TvV�%�*XY�]��6��@mv��M��0��S*H_ݰ	���@�fo�)cY�0ⴌׄ}>�2��-a�N�Q�.S��z�	GL�R�*�sJ������<|Sh���6+M�T;��T�_ۋP�Ί�u�1����ɟ�jK~Y���^��G��>ܖ,nD&�!�_��2Z���TO��ȼL�:�-� f��]4Q�FX����������TK���ӭ��?gnЖb�^ŷd�����j�����kwrc�S�~�I	�ZL��dK<:83G�*m:�e_Ğ�`L/�m0��5j��Y�� N�
�CC��Knn�,��(�aϑ������Z��f���]��BG��5\��;z�܇<���y�z�j^����ʉ�Y|�Hu��i化��L�"u�	����>e�e����3�<����F9&��G��U����hBJo��)`�rE�>86Qb�{���ȨMMF������B}0���"���9���"�p���0�:q�BM�r�6�?~�y��ߡ�̌j�*���N���}���E��{��es���7���'8sivyp����o���{ta�:n��ю�5j �Ǣ�ɅM�Tf�D��iM�F'u\�#���Oܻ ��r�_������E�����/�����<���?��798�QO��;kZS��R����톻�"��3���<��>ʜ��ΖK�-����e
Z�%^���N��A����w�|si�=��t5]���l]<+�����ڧO(,��HĻ1Oa���G�c�/d�8����B���.�D����%�����X�_r��g�b3˥h��w��Y��۶5�ʧO�,[j=d��C���HyU�����i2a6+b�@���'��э�E��_JKw�*��BC��#����Ɔ���7E7�:�]����b�ym�!jXo{�ƟQ�i�R������چ�;Bܞ5WZ��w�*t�
=�P�z'p�bm��N��^aW�S��!3#�T[?�!�n�~^�Wݏl2���<�4�M�s��r ��<�/��=�)�>"�Q\эf�������76��GsX�A5�.Y�n��Gi÷��q����h1������m���)t��0���7j�L�|4uHɬ�p���<��\q�+.���[y��#	eϞ�æ3���~n+pN�>�N����J�S�4�[�w��Uʁ�K�aG+�Z�91��C{s�'�iמ�:i��A�Ʀ�������4��*�:����:KTԏS�����������K*9P��CX������G�Y?�m~�'��'Ծ �<r��;p�^��}�d#k!3�Z�ڝn��n�?k���A���>��@[�����"����5F���z)��޽(���_�}i6X�~�����(�m��`1xq�ۉ�3�A6�,���"eo��:9;!t����ם��Ǯ �pÅ����V ��rx�'q���ֺ��,J�X�)1x�k(�P^��h�B�c:q�C��u���A���p8If"e����P�%qJ�֕�໧��"���ɭ}�3t�4<�>�ac1�o�����_�|+��jp�%�z]��@�J45Qq�#@�>c`��r�Q4����.����$���yv�-�4�IUJ�.���Ѯ�8���:��(�ЇuWcky�g��I'��?ܴoLѐ�bA�p��f�6�m$�bxk�06�va�c�ħ�7:�UG8�v��)J]G�OY.t�vT�^��l\�G���a�������^ckq�����_��e���ǎ���Nx�%4���mn�ty$��.�f���Ӟt�mv����̠5l/3�w��O{��b�O�������{��F$�+�?,���˖��|r;�R�	����dO��&�Ǐ��zה�V��<�J�[(���ɼ�a�-��1�O4�9��&3��n��|Xm+���;������=�ia�i'e����ym[���qu�wV���@51W��u��GS����\>%�s_?Qq9o��BZ��Q<	e8+?�0����[���ﯱq
���-�%��c�{u�J��sF��Xt T��O=S0h�MĦ�4aWcc5Ә vw��������g1	��¬�*��mS�x!�����S��!�HVg~-^o�	�/������_8�|g�O��5 ֯^c����|u�c7 \a�e�5�%.)�����hvB�o���*c*|���l���o�reE�4$R��y�������ݾ��%�#�f�W56������`�M�y"D�Ž�'N���̊G|���P�������^ _93��S�dBh�¯�=Ӈ��
����W};��.�<�ix9�s��s�3�ࡏ펞;Qɯ�ِ��4Z2�G��~5�PEھ�Ҷ8�3����#��UZ~g�v�+�<�����YݒW9�`pn�b��l͔���\��M����$�<�`/�I!�T�dP���0T�gΊ�u�^��ʿ���/�Blݍ�������݈0#0O,8��l�~�
-�[T�[O�_�'Y�Б�r=���7�᩸�`>4	�����`�f�,�W���Ħu�3�0N&�Ȱ���?w��!�*���O�����.�*�`%�pUw���ڢL�Q+��?���*�H�y"ײ�n_O�r��??J���Q�|��a }�q�C8yk���k��A����$�8�[�]̩����Ѫ���Χp��ZfF�l�0>�Ϋ?��-��f}��o#��}���i��N�{$E$��C�AUh�M�Fe}��o��o#Vwz��U�{����&����\�w�sk��ёo���Z�R/xJr���w��ԟ�%z��m=�t\a�1���V���
���5�E������K#�f�/-�i~���!����+I�#��;�O��=�xEU_��������W��,�!�1�S�vP�J��t*�_�X_t��e��m�r��+L<�L�8�y�X�i�7�U=�.��ԫAӿ����Y�³f�ۮ�n^��Ɵ�ŝ����~K�?b�J+�Q.x�i_���1ZLM���m��U���K��@�굶^C8��:8���č����*K��SMǉ�K.�����*D.i��ˌV�y�q��\�*����n�C�t<�b��6��3'85���~,61WQ�ܕ6yR��P�C׀q�'�'�]�--�Ứ�b�j���?�U*��GA�'Ю%�����W�$;��ϳb�u4_s+���!�1^�Dst�ujr�V��݈��`�=���/��G)�:Bo�����Z`�q���zk%��2MK���u�0�\z�ǘ��u��% Ý�[S��|qB���|`{�P�mv4�V�G��g �[9���e�C�p�����P����=�3����@��,���$�3E�TݦZ?΋M�RC�-y��K��Ok.F5�����̗��?�OL���\H���}��~�55(#q���^_rJ� �U߬��uZ�cDM�c�5��t�.##���-�@jr	w��8E�g��9��؀2�_�G�+�O��ncrZi��
�5Vn�f��;Z�򋫯F�@��Fq2���mO��RY��C]���p����k���T-�H=�XR|�Sf��G��� ,c�68p�B����T~.P�cUr�Ԡ���ܟY|��W�V�Y�ӱ@��q�ʕ�l���z���\8���RnK�?k9�I:�.���W�C�+�����˄��W�,z#2����N��;��7��)[��__y���k��FA����b�������}�7R�O�8�>�Fa4=���zo�J�	�]�(���'�ޠ�M�pb���/�!	�����0؟R?�����j�!hhq��4��&�[brp�}Ɛ`�O� �0�L#�d5b�clS�P�V کYZ�\�6:��ȿJᲛZk���ډ,�*�+�.�gy��S
dw2o���Z�n����XA�eބ�K����Kƥ@���z��2��7�Y���
e~����>�����?�����o�0�"��!ic&���|IU�������:��o��2��=�H2
h�"Q�b���<�����d��S(8��0�s낽*{J{�q=K���џ5MF]�m�)&�(��AbU�TR���n��]7�j�����qI��
K�-���ۙ��ên	O����0�+:>7�KbF�SU�O������ȱ�uw���%#��[v*��/���DW��%�oWQT���/��Ш���LJ	�r�!0����H�X�ϯ)&���|��Kq��n�?��zȁ&H˳v����/�\��	D��_й$���S�u��Fͼ��7��H�u�t��s��2,���j�}��\��k�A`�./����V�:�
f��\�7���9��	��3����C�^w�������V�����xl&�c4��#�w��}8 g��{���sz9uI���zD����y6�cWR�C�GFff|�����4g���ޟ�	�#�>%a��o�TO����<ژ�n��9d��v�m,[�m�*v�H��3��1���e+���.���"�T��?K ֺ�����c�+P��"��H|���ȃu��KY��ML��8�L8�A�<�[�{w�S�l"b�g���J�I�z��O���M#���*��2znx��?�V�p�:4~*��� +o`e�h���~�81	�F�5=��,@\�ҺG3��'_%�'�'b(�@�)�J�Lx�����]�=����v�͒9�"�&�5��i�z�n{��1��v.r�V0�6`�x����o��c����[�v��c�O��C�c����\�6� �M��!9I��U��N�	�E�N�)Y�[�Τ�K7�4���K˛߅��%���C�Ș���b���+��Z`�lm���9 c���vt��kw+k.���98 ��eyIɤ���kYY`)�Ȫ�a7�����W;ڵkυJy?B�".eœT�1C�����E�����������^o ����WÍ��l�k��Y�Ͳ�_+'WR�O"�N2���Hp�[��an���G{��V�K��s�E6�M)<K�P��f�߰ tqC��=/D(�뻠w�n ��6�o��� ��*O����^T�Qsˊ��=���ھx��-��/�gA�rH�k�$y��}R\��UJ�~��|�' �ƪF-�Ƃ�AFѲ�nEՌ���?^z��t^��2+�V��s{E	��+�c�#L
l籬̔���e�?iK�N׸޵��ؠΦ��J��Θ�!��OV�؟tR8�`�E��'�q���%��Gɬ���:��S{��e/��'4�<�֢��"{䵉-g��V��,y2�sa��ׁ��M&�3\�g3S��Α�5�c��?�ۿ!�C��d��R9�n��u��G�d�gd��̭���/�fdf�P����U�4�$����C��/�8�Lp}���l&&&�%Jp���7�3�@�Q�I��N�$r:��n�.��{����	曶�#�7�q�fg�l/^"����/ m�Î�y�L'�B�D�/�[�cF�z;)��{Tii�.6�f�m���hÞv�-�h2�����
��Y"Q�����(���}�c�HO���$ ����X���Lr��PV�w���j��hH� ��,�#�r�Nk`�R�=-u��f�^ԯ_��A�xz7�N���q����k��پA��Lt��=�[����]9@W|�G��ىQMNҿ|�}x�| �5ie�v�r3�[M����"8v��^���~��p�6���y=9g�h�v���`j�]6���	"˓��u�d��_�G�͏۟���7U�0�n;���dY��wiȸ�+k ��y������=4.��1��x=ڽ�_w
�b�;�פ���C���m���e@l�w�*v>���I�~�� �N�ݿ�;�7�0.�}��<�֥��>����ޑ��$��6�����P�B���&���kC�3Aa��X!�b�$ʀ������M۽?�I���ϧ@��>�5$W�>��P&(�Ŵ�B���=�	�@B�-�U3���h�b[�4�)(u����;K���-#�I5/�,��(�C{+M﷞�	w���&�	^��wq�G]U��cj4M`׺�ߕ0�x�}A�j�\bŴ���<HH��6ݭ^�L�9��v��PZR��	[5@ EU�2���j]2gZ���`K3��Z�c��bK�.gY[��w����|�7�]�9�==��*ItD����t�5.Is�P���w���5Kfsx�ķ�]�$��?(u(��ȓ����^�z��@N|^UD[��4�C4�i�ɏbpר�S HV�x������a��	ɸ���c�)u��+.���?j��έ��>�x�ؾ0o��7vAC�D-��t�X�I�*�:}�[�U�H��g�o���f4,�����׏.�ӗ<�Q/KwEG@?��Z�t�SU�t2]�t�p��$�v�1U���~ɯ��i��Z�Ѡ�|f"8�
e�\c�)y}B����$0�Z���BQ�!��X�D3�Ȃ�G{]�X�LL0�Y�'���(X�tFG�1�[��l���2
'�%[6���I��7�������-:�M�g�c3`1=�n�:�54��:mޤ�`�y�Ǭ������E�:ߵa9Ucҟ��w���^p����=����N�X��\�/���N�H9�l�f8�c�0�]�����thdl{����RTWO,�]��A��~������"���i;P��t�k���kZ�,V��0��ʅs���z��YtoWaȫºޓ��˓�Ę�R�7�m�g9D�����{V!�%���0}�
�JuFf���� �7��m��J��L���ܰ�Z-�I��]̆�V�tf�������]���X��r����74��na��BnU��\5��;CTR�cc�p��� �n�3�� �G���?��~���Q�ι��ȖZ�w})����vBD��{���'2�5�&Q*��'�S�������M�*�Zr7����_�%�V�T����NVK�,^֏����Q���Ȯ��Ɉ8;�xZ*1�=�Б]K��4�n��Z	V�1��Rs�g��������O�=q�����d��dܟ5o�m�U�^ur�#U��Y�>�<�6�m��[��o_�޵td�� [y掴ʤ�f���$F���U�,�-�K	����ȟ�u���3G����>�����<�2�bu����sWf�r��r��t�f�`@o#dK���견j�Rq)���4�/�S�瑁v�eځ����fB����*�.�6V;�#��/��Փ���嗊�*�H�Fh����%�M7��=Z^S=��J�k�ȉ�K�r��hK�%O5�o��;*S�6u����Y�����y�*�������S�b�q�n���X���/�imRK�0La����մ$Y/��@5���.��Ex��)_ŋe�9�z�1֧ђ{w3$J�E\�0��cG4vO�������w�w��o	����s����@R�}�K�[]�Po~�)	�S�j�ݗ��m�I��21�#��?r��`r,���-�z�id���q�n;Ό�iJ��}�6��8�X���@w��=Y�`OY
Zw��y$���D)����?I��\�UP7�u�mIa���l*T{�s&��2��Wu������ȦKt�Yހfl�I�*p�b3�5vb���-^m�ؑ�̢����i��ȼ���.-�ZA�:d$%��9���T�ͫUA��"���Z/�5�I��;{��5�����Lz��G���4�Um���׍��O ӣ�
�
Sn4��g�q�N���R���7�K�(��,
�ڋD���ղe��⹶���_H'��fl��9rף@��mtT{��܏��˻`Ɵ9{y�/Q�ti���LhP83��_�
e�Ae!��p�����oXe��66��9(7�,8��A�Ճ�Б���Pj�{$�C�������~�NQbf�y����� X[���xwP�,�K.wa��l/`B��`q^�W�Km^�O!^�U�AV���lE��-t��cWq�rZ+�#k����V���Z�T�V�!M5!�����[\SzY�����[_h�?7r�%�ϯyۄ�n�0<��3lKSx�<�;��~����4�6���-�v�AVcZ-hc�)��cb#k�0#���1�ۄ(�I�kދK�I��/��]��C�q6cʞ_ͼw���R��(����=����LOR���M���F-A��M0F�ҟ��a�*���mbϟ�2�t�����;�E�2�8��p��|K��zq�&Y*%�?�ߴ5*�����֕���ï{�2�S���/�z���$cG��'���?:u��	O����ՊمK��u��8>L��h���:!��=��s�7�9;|�z쪺.�0������HV�����c/k;<H���T�����g	�� A;08���-O�?���>��{�0�u�	&�Tq���Nv������t=fmkXRU��۫*�
}o��3�`'���RY�C��қϏ��|�p�!n2vSп)�;flL�����[}�[,�YҴ���i~C`<�GȣVͧm�پ�����/�gjt3��NX`2硊��ͧ���v����5$o��sg�ԝ:H/�J�]N�m��8�����h9|��o�LWB���O�tn�h��:E�0�� ��Gg=o�n�ǖf�>~������ϲ�WՋ�֭�I̷x��@7�[�r�f�1K�rq�Y1;����5S��P�F-�y�e���۫s���$�o��`N#�������{n� X�c^DB1����C����g���}_kOs�����b�mT,sg�&^T�6 ƌ�*z:��ݪ�(�����������U���,�i�K}���.X_�of+O���cO�7'�h�{ĝy@͞O���Se7k�T�"�b25W�X(i:p��Vա��z���ɣ��I�}_����)V¤���e��ysp��0QAML���0T���o�wrK��~Z��i�`;�MO脸}�ች�V
}=)KE ��MيfwQ� qN�0���*X���9���]�d}"��9�>�H�\��Oc\}_�}�'v�-��b�&N�UL�E�R�G2��lb��<d	��J�����;��i8�9j�$k��Ѝ���B�?��$��2H15���#FG��k�P�<�y8W��T�i�l��0�b�i�93��4Yu�pϙ�Q~W�!S�9р�����7�3�]���$��P�9:�h��P��.r��8皻?�0�I��E��ocl��з�V
���1#�D�;~�P�൵c����K�.|�ϟK�/�iu�5��kk�'��9J^��	y;å;.g�d k���k���I�wT��'D��~�]U\�ՙ�(v��_�}�	�|�����XfS�Ǘ9q�1��D�Te/�;e~kb����������MA�J0:���t��2�1A�{���>G`��� -�D9�3w��>|1B/<�z�L��L ⓟS���7�a1�ɓM��
��֧��k����q&��?���:���Ji������s�,@||�p�s��������s�e��	ۚ[�����^�e��a�dW���қ�Gwz�����E���|���!��*��!�a�h��j���IN�v]P�gX��ml��&�u����hm�3U���h�6���@eWoy� �Z���7��Z����u���R�1�q���3��~�݂��������7"@$�Vc�(��A�礴&��!�m��B1�;7�}��>Y�P�f$2T"M���k�m;�vPȯ����Z%��󬱒ח�\��x���^%K�\?W�u��v��zD����
Ƽ'�	)aZ�C���w-ER6XR���Q_ �Y"t���GɅ��qӹ�;��0ݥ S0���5�P[N� *���a1�eF\� \���6;B��W_�Oa&P�m�XD�
��$xj�W׭E�;������N[��E�{���pǶ5�@�g3,Ӿ>�^;5�DGЬB��H�Z>A�x
������}�5�����U�X���~���=jfZ����:G�jX9��	�V����t�ң�] �l	�a�x*�,
^=a_-���@
S����i�n����H�]��l����!�BD�Vɓ'� ��U4np��f0�-��i*K�5Xv�	�h�</�o�c�x_�kLйfWò��J���U\�h�I��U������(*�a���TL�#~��B�b7�)Cz�_��h�2�����|>Ɛ-�}-�G�DYn�͟+B�y��'�p`�cp�F�_g�R��WtBN�8Vp�G���S���:�>:e�.Mx��-�M�E�ڲk�V���cm���շ��\�	�EA#ȑ_��O۸1�A���V>"��	/p0�X��J�K)ɯêc�3S\�ոb�iG��W���g�ϲ[��3���s�D�3��d��Ϟ�TC�RI	���Y{�]V�H����i�7+M�����-�a�J���{9/&�cJ�ԿL���>OTm��o��b}�WlV�D�f���C�����p\�ӓ Ŕ��m�JuoFJ=�����;ױ�ח�8h��:�	Qm�\/"����N�8��g�LH�����/�)@GIU���Tsq[wξz�v���P�!6k��,��]��W�_6@�9M�Cw9A
�(��ӓ�����ɵ������Z$�/�^�@5�EwU���B���=���>
�.NePm�*ǟɝE7��Km���C�c0C��n�8e�����}5�v����V���0)۵��4��pm����|�W�8S�����9uIJ�fc�+;�0��9P�N6�"v��x�U��rz�<�v�h�+�_%VQ�T��{x��d�0�5��/�_��U^}����g��~G}��D�*��q��;:*������LJ���wA��[����D~'|'|'��!�r���^���>JH'�����7]<u>ԩw���x���w�����d��τ��������f{�����k���3���;���3���;���#X�	@F1�&BR�L�xukk��&5! ��֏��ډZے��0gŌ�r�.ܝ�����~}���ESC���s��C�G��W�~�}�� PK   �	DXP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   �	DX/0�m  `  /   images/f42dd85b-579e-4617-aa27-44ea24c5d2de.png�yeP@�&�H��w��]��!����}qw��NX܂K��x߫���u�T�t����twu=�LG�(I���������H��k�w�C�ϣB��w��$��
C�����P_$t��qSw�t�4u�����d�q�s�j�d���b�u!HC|.+!��}n�@���ftw��[�dk�}� �����J@LMA ��s	�s9p��%���Oz����P��&��``��)��<6����!9F���j��܋�Kߍ���n�Fqg�Y�j�Q�k����,	d<�� ��XX%��PB���&;�<� �C�B��}�D3�#<<(�&0�ߚ�Rq�2�H>7�x�?!���6�5��<x?j)�!�YP$T�Ҏ٩&#͂N!��lS���T�^)Nt�헳e�p@�^��[�S[`��������|e�#�A�gY�n���<��h��N��.��)�ʝ��.���A�lw/�\ʗ|بp��V���1�ߞ9���ТJ?)Z"8���<���&�@��J����P!���w/�60�լ!fI�v��+p;���mn��=���Q����z��i:���b/LB�ӓ1CP�UT�
(���b��(Ɇ��������T6Jp��=]�����$�N�u�A�dX����]7̵�R�:��c�;iV�@�!��B������x����k����(B�c�,I����?{���׉�7�C;`�C�O3��/��G�/K\�X�B�Fc3�	�f1�A�aj5b�dL�a�嘢qxď����'<W��b,I&>��SעK�0�N��e|�6�_ �gm���~;;;Vo��S��G�^�ߔ�G�=}�U��љ��J��hT�1C�{�0���C�&fa&2^�A�" g�/��C[l�p
Y���R�F��lR�.��,�� �	Na">?�7�q��Ճ'3�u�O�r�/��^f=9�,�F�s�^ǧ5���h����s�_W����@~�n{�q�\Ȅ!�'RS��4+mk��ͷ��^��zx~+F0��
�C�F����E|rz!�l8fE��Ja���~"�����q)t�Ŵ��O8%�Ŧ�2�b��>��8E2���[7GG{¢(A4ɪe��P˪�-#@ �	�A���:D�T72�x�>�d��&Y��2}`c�!����lXa��Y����e��� &i�	:�J��{h��;CO}�~+F�7�����yr4������WG!�3�_�D���+F9rѯ���βh|E���4�ޟ������v���#����g~%���n��Գ�j�����W���s��pa�֥<L�Im#>Ĳ����)�@��5u
��������{A9W�M�DmnO��<���5��Ā	_�o�zt5s�E�F�s+�wx���c~�]��ǐpJ�{/yڡ�Þ��R�?SՆ���Z6���I�B���R�LF"�Mbt��)y1��F�1=B�(�R����/=���T9gU�R���^1�mR|}�Ƣ�/'05�Ie&�;l��)�k��/lP(��^�Nq��Ca	���c�g�Y{�PSS�t���#ok��T@��H턴X2�b��66���bKGvW�)%@rJ��--�׿^��[rl�	�VcLU��%����.���m^��{���C+8UH��_XA���Q���9q!I�����;z��߃����]��aa%崛!Uz����ˍN`-��S͚�*����l��M� F�-dė0�&�Ljd�I8�!�L�C2b�Ȯ�޽}E��/�}�?���'�Q;��k��k���;��Ms�4#ꓔie'�s����/e���ȸ%�o���}Z-A��KcO'��)ö�����fT|��������<+���N��9_���/��3g�(�qX���5�5��!E��]l���g�[^򀉪/!p�Ȱ{��,�CY
�=�[Y2U>R���i:&@C����[�*v�+'����T��t��MҜ���H�����`�W��Oe�de1�w�m�З��Vf:��g������:�5!v�,vX�"�[�)�:h-��k*��+X>����o���x�h'c�/,Ϣ����E��?j�C�e�1��򯖹8I�|X*���6�	yD��R#��%��7f��y/ø~�K�2�;��g�R}>*��i�S�Q�sHƳ�d��.��h7@��֤�Xw���bFQ�����$\�GQ۴��P��d���Ϩ�'�7�Z�����msZ���O�~��{x�ܙ��Tw�ոS��c�(hNn�N�-��6�(2:cf��qmpQ��>]�Q�М�]��(jZ]�"0���$�"CI���&���Wt�W{��"���7]ڳ�&'�(��
�6��KU�4E���g����f�W�.6.�:���d��,_\�,�X^��A�\�_��PZ��,��j���A�~Ejk͎��q�`��C,^1��w�F�?���w˺�Z�����u �h�~q��ZͲä�<ʮO_���c�R,�+�+��ٳ4�Ֆo�T���.���z���(@�GU^_���
�1E�����;����W�nr�N�G����	���X��	2@	1��f�I*�?�;�a�q�ܘ�����,�!5���C�d�_ڮ��x�~7$�=�ήf\�����&�l!D.+E�I�k����z�\*���x��S�1�i>����T�W��!8�g�ɻ�4e,>g�=����_S�d+�i9�w�a'�?�%��q���k��2��0��YK
v~V��Ll���Tx�L���iKx�&�q�R�#�_A�ߺ͊J*�ݼ0��/�����43�����1��t���<�b���K��
n��\:������x�\�B(��z�$��F{�l ÂgR��7Gޯ[�R0R�u�l��T���J'���r ��3l0.�b��}]�3Ѻ�8Ls��jAvl���g��s�qH������9�{�.��4ި��!�V⃪ߞ��嗓��¦��8�`�h�1x��8��'8DM9z�]��$MI!!�5v��&�I�2���]j
��O�FFEd���$R�Oद�ټ/�Mw$��X�u����ڬd2��b��Dՠp�TK��;&��Ω�~rl�#R��WS	��^i��]��A���;|a�퀽�<B�_,��_d~��u�v�03��A9��Y zY;^��Ob�� ��=x���Nr �yI�b��mG+����\�;��=2:<j8�[~8�]n$����T�����!:v�	{?@�;hG[fj�ͻ������o�YJ8�p���|�i�=L����|)Uq#Z�z� I���T�`�K.��x�5��y��5�s0`��HJ^ȉ�)���ݲ_<S	.ӵ�"���;������1�&O�R�5� {k�g�sr1��;	�tE\/�LsK+X�� ��i��U��;�.��0L$U��p#�GfQs��,���U�����y;Z�t�>V���	3��x� ��|�Z���RM:Y��|t�h��>�F�$u�S#s\|`��9���y#A����^�W��$]�`�o�"�(>}j�+�bԾL��ו6^e��5n��̷����ѐ����_E��l�J�}ؚ#o��R��uv�;'�{;]�.���y�P�L薤n�-�axS���)���&� ����;��CP���	G]}�ձ��;�]6J��7;�8r���π��q��O���ٞ=Z08}�z��I9�����a��+�����-.)Za��s)�͍�q�稧2���;t�I$���b����.\BW#4Њ�m�6����]Gg������{�=��7�H"�M3c*]���H���I�R���"�T��j:�!�yga^2����)ñ�C	�#	��x#z����^�G��[/>��F�����l`�Ы���/uLE�f��X��;�����)�QY~��?~�k�l�m�I��$j@-�ڐz� T+��31Z��Aaݗ1r�����-$^n��G_F��md2ø(t�r��-R���&��wl��I*=2���N}]��Y��~�N'b��oɕB�'b���ʖo��'4A�'�[��ވ��w�Sj�FxsC\f;=�[cNA	"=W�@z>;7���� �vѺk��W����w��0��B����@�u\�hٜ��3���Z���p���%���V��G(���h"��Ȏ�1���X�l�����g�쾠��:��T����=AWܐ�=��x�C$�Қ �&�%�͠�<�Q�e��n* �o_���{�����>z�p��0��w���6��81B�v����ʮ�/��o��;͇�n±i|�/�6����סiL�伋κ!H������g��(�9[7�6R�*�D1ku�Iw��l:�Ĳ�5��iJ{8�s��Y�a�WF�	�C�8�dGc�.��A\�ߞQ�~7��l�t�Z~Ϲ*6־��&������\�j�~
�cpC�U�og�uW^ƻ�Fr��	dK�D��,�f�%�`��[b+S�k�E�ۥ26��,=\k��P� �l�����A�V�s(9��\�p�v�=���/�ֻt�d��H�wVDw�+���j��Y(�M��~��+����cv��͙�)�z7l:�ӛ#PL�B����l�0���pE	���&#�����k�< h�{/��Pc*�x����p�/�����;"+�)�.��u�!��hQ���c�A����ȽdS�A���'��|�+�}�@`�i��! ��|�6�^���#�G��[��AI�L�L�������b��Z6fa�d�_�=k�9�q�s&fp%њ<~��9.������Dr�b*�O�) ���	�*LH�p�-�s��,͓y,`��ж�sR���"	L�R<�Z�Rɡ��	�*:d �T���P�d>�� �=$��kwGږE�upz7TM7��޸J�� �2>�@�	��� AgX:4�m7�<P�t�i}P��5�$��
��LMtY�я�7'�	)#}��{4�f �3�������A�9l�����MR��?'��Z�s�Wf�FǺ9����Ld�j��\��ƪ�Tc��f-uW`�ѡ���e9��t�ƓS�aK�
�}�.�7�a���}*U��jy������S�#9�S�>�DEҟc� A_�o'�gm�������dR��c���_��V���O�`,�]K��%��_~8n�6���H�4�M)�� �?n��U����:�j{�<��GQ滉���koP���v+j��#[>�����!�t�n±�+̺<�ታdKGJ�]4���nG=��D��{���
�k<�z�����Z�S'{3��?s.������XE�9���:%�}ڃLd��KUw�����4���[�:����]ŗ.�jq����/.����[!�,z��Q�߱��B�Gr�Z�*B����`�ۘ�|=�}�Q`.�$�&��Z�v��䢕��!{,;Z�A�ȯꠕ�O����3q��;	j�R��\�W�n��*g�'#_ �8�a���h��l�V,|&_I���#�;�D�<�4W���u�=T�|��λ���|#��u�3��t���"�8e��Yq`x�h�}V���.���zA�>��ŗ��8�y~]�8�p���S�I���ߏ�#�S��.����W��1���N�����%�0����=V@=�:L0��ZGl�Ⱦ()���`YS諯�U3�)���2ʠYt�#{ۂ7�`��?h�Mn�gioi���(�#�дJb��f�˓�ln~��ƫ��&~�xi(�o��<~���>TK�L��c&��œ��aG�k��TR1�s�j����B�ƽ�^R%�x�_CK/�r�}�?����oQi��Bf7���(��U5��i�L�R����k�����_����X�W�Y��b� KFS��$�U��<�-ƒ��X�_�BJ�o��;m  �B&�gM��r[�9�f{��T\3�i�99^�:�sL��j�qi?N/B���
�c��'�D5����xG�x�zt )��֑�^�p�;�ݧIS5[�o0ǵ@�x��m"��H5��[Р�gN~dw@Ҏ/N��lu�9F�*�^�GF������]��P��0Яa{��u�;ɫ�5��/���4��m	'/5g!���V:���[�����������)<4�K����ƯXSn���B�����*�4|�+l��E�2�9ڵ�����i ��#�j�dD1�YIz-{�7so��:��'�����p��`d^7�#}���"�e����ci��ｵ����l�ק֣�
<;ϻ������o������1[��.8�4��->�!I�ܙ;>DHY֋%�:8wM��@WtRR��?�?�nW�}on&�ȍ1�桭�q����/ۍқ�������nLeO	��>�ݼ���W�)ӧ���� �/	���F�eG�F3�%V������i�]i��]�y�n�A��0�^"����_��װ�3W{j�4;�#��	� �4w�[k�$~	��'�1S�M���xu9�X�M¡�5ZEr-C�g�c7���u���z�hn�0��~��K?�wcL�P����hv��b������n�N�&{��H����ӷ�C��ݚާZKײ���i-2Wc��y�,j�������y���e9{RS�p9K�=��N����5�ƂZ/P�C��7?�v�C�I��)/aU��i7��|����^�s��DD���=���9�D����ո��YTg3�E�oU&g(��T�y��:!���V2��tq�����v�z�^��y"%"����pڷ�q��ad���:�a���YM7ŗ��K��'s�:�@�����G��y�xj������t����l`E����*�؅����q��V�Eт�9���^2� �[7���>��������y�d��	 *�'Bpi_���g49�멇��H�"GE���J��L��״��߁
��8Lkn�
m?R��[O�Թ�ԡr+�_�J�[p�Ԋ�F���Җ�M0���`��Y��-k��.+�	���S�����X�3üYI%�1���PK   �	DXF���?� Q� /   images/f590943e-678c-44eb-a174-3243ba5f3820.pngl|	<Tk���ܴ*�})�F)�2�t�d�2�L������'�m�si,Y��kBc�Pѐe�C��4&��4���ֽ��}���u�s��[����9�~�і��!��sdS%"�^��I�J�<��}���z�߽�7���7x��BC ����V5:_6(�ex����������__�C�n(��u�C�w�Rg�d!��c�?/��}Ƥ�X�P�#�}�`bVO-NX>��)��l��T�z?Jo���c�!P����[zl����e�Kyĥ��j�������v(~9�9�D�FWo5�`�~NA�L�L�4�M���-;:�6RT��!f�Y� "��!ɱ�����?�snRr�D��n:��8���0Y�T�Ip��Ҝ�Q�A�-f.u<��}��Ha9�:�C#J?~��X��s&�D�W��t|�ljt�X�g���x<�K_�C�LV�},�2�����Yw�揹ճ�<	WF�x��C4[K�9�p��8�愝���c������4r�3�v�R����X����i`O���-��LȊ���G��	H������hhiu�r�ׯ_37lےlY���~�Z4d�6�I�革��)%�ͩ�Q�[MF�)�OV��n0��X3<S�/}K�M�8hD�2Ϟ��s������ ����~G
+���i�j�[ZZ�c�cta���{ZJ֡.�����m��cɵG?�Zpm���k�����9ׯ>q��U�X�Y�P���Y����_P5��a*���z�$LT偽��;4Hè�<H�(�?�t2��s��;f�9w�O!U7��b�+]�){1K� ��"[]�c�d�z�0Oa�[����s�>���2(�|�z��[�?�����
K�9n���&�J�����Q:���rrrF�
�^�0y���ݾ��P�8�is/3���CE\b�m�7��'���%젡A�֝��)n�;o$�)Y�?cd4�����ǲ�W���4�+���H�V8J�&55�iek��	-iӥ��PW��*��CCz~�G_7Źn�s�_w��G�m��ϋ~�U�dkih�KjC�]1� ̈W��0�펻�Mx��������$M���-L���{�����u�B>�~�Z��"T�>11�+�������В��8���B����l�C�:4���y�;�W�$#<�$�����S�z~�"2i>5v���Є����� =���h�[߄ɓQ(��	�o}��*Q�=�9�"�V���� �*�6�^�V��k����:LY�Pc31�qP,�«�gZ�����V�vЈ��$�1؂�|�]4z�`'�mB�w�F=��[vo��0�����\�����@������m�W����ю�g|S���q��f?��p��5 3C�_��+�'�R�?���Y�S����GLE�����	Ӡw��qa�d..�\�z;�m�:==m�����4)g*�*1�d�a��������'�-F\�	[����;����k����!�,l|t��b^�z�����*��+[w�ҕ��Slg����	c���or����Z�$�*
��@�����mq��jPG��5 ������K��}��v��q�X�=a7Ƀ���g���C�>k�Mi[������z���$���wk�Υ䌔�|�����Q��w���9S�z
79�8W��7�<����ٗ�fh7kM���0��X�>���3҂�<�B)��֋ZK��uF>&�<�2-hjjZ�|��T����-�2���!�xF���K4즕O8:&|Yp���S�{j�2���t�J�0�'���5�ZwX>��_�/P��3;t7��co�ȉ�Ŝ1��C#T��I��N-����k(�KR�
�:y�q��9�N!�.?���s� ��j��L�b9��&����?b���*d�C4�ew�nU`$aAE�x�n��2e�J4%!�d�.������8	�MCVBP�!���f�U��#�g)�s�]: ��������chu�u�(#X�R�h��M	�%�Ȭ��HE���J�٤<�,�#��B(Uc�̗mo�r!(��	�'�s��I���`��BBQ�K�[GS�dՍ�
(�C�ְ�n��m�n;4�JZ���|٢��i�]V"�':��-�����|K�s@��'��` ٿ�A�k
��~��^
+[RJ*���c� ks�vxpQL�� ����&��4"��Lb�%���	��w�`��i�r��
��"S����-hw�5
��B� �x��՘�b薞��;�(_8�\z��z7 �\����u];#�U#�ΊYY���Oꅄ]�������N�n�.]�!k�ϤZY3�@X��ϰ*9�	���Z9%wd-��m�C[;�Vi	��gR9��YX��1AŘr2�k����I�e�oL�c�c X�� �$��I�-Q��3��`8	YP�UsA��O/o�)hn��]����H��y�H*沠���G�F�'�b�U�<HýN��z�{y�ʕ�/kk���.U�iC��N�e���lmm�}H:L�W�jF����I��u|�OB�*�%g	\N�m��vL�e�Ӷ��I�A�4�����_L/C�I�h�9F���*56�!�UyO,Uc�P�r&MQ�e��5��s�TM�AAW����w�+=�ב�5�I�>UNva���v���������%:2ק;t�$1yX��w'�7��9dڥ������,��ij���dV��?�*Q�B���`�3~#�	�/�#I5AE=.#�}�W!f'a�9���Y����~w�"(_K���Q��
�
햘��2{ s�M-x�.X���%R�NN`Q��,�Ȭ���%�K�U�xʣ{����o�?|�y���Y���Xe��ή���a�3�P�|:)_�T�8:�<�����%VUa�����ci�������ɒ^��ީHP.��=��WJ�����,w�()��
HWu�c�&d�=Z�ܢ��V���~�
g�HR�����J�u(���5����#Y�*��V����g�����h-�4�͛7�C�x��m��w
����^����~��Et�̉�A�P𷾒�T��״��)~ޚ~�7ԃף�W΂��HU�����\`�ϸ�Z�s:��Y4]p��H���q�o			�Qw���q�� د�`u���O~d��2���hJ}�x_x��V*��xcE�O� m-����f��1��\z�[�a���5~���q��
�~���7W��i͚#?���t[�74|q�ҴO�~--U��~�t@Q�5�5J�^�Ч�%���A�Z\Π2�[l0Ӫ���d�_��ͥ[T?/{�CXy��d:>U�-	l�"[)w�#�Ȕ�4\&�Zv��GJ��>ё�Z94�7�ݯhJ3���$O���m꟡�K�$�Q_��Rą&$�R�U;�$vu*���Sæ�g\,������,G�.����ڵ1�S��T-��K��j�#\�����]-�E?�E��a8��C��N�[1�ND&k��M�R-���ʺ^1� R�\)������oʂF  �W�1Z�����Q쨿i�P N3�S8%a*��L�f_r~V�b�+��^��G�PO[ͬ�W�k^�0��:{�R�^�?�iW��,���&�ciG0h���2N%|K���h4���{>4�Җt��C  �L�u�uu{<p�@1H\�U���_7�V�������A���w #��z�Rw��T�KR,έ3s|f�!I�_ܓO	��֥D�$YY3������41�}��OCכV���I"�a8# �G@���,�~]�:�<Y�f��ے|H��R��a.�Ӽ������TA����MK�u"9i���	CD�W��~>e���_v:�v)4�4"�'%x���CG<[E��������圲�m�»K�=���#�$ǥ`n�?�P�O��K��m���Zch��m�̅}�����U1O�"����8���.�X��/s�>����&���50R���V�ڏI�pR�&�Ӯ�y�Zk|��#U��I!�^x�f�pEo��"�!��P��@�f"ml�&�v�릓"�%��"����JZfv+�AO� ���2�a5^-W�K�C	bѝ'���.����Z�r��/ՏرI�u��&��/Țī�d��s��< x�B~�����I=j��dA#0$����Ǥ���P�)�X3���Q�����i�z��?(�u�9M΀ѩ�@M���j�#!��-��G&�dD��5S!U��s��C�$t̘�i�Q��w�_�����1W2 ��\�V@�3�f鹱R����)A���;���p�L~d��(?��%�Չ����G�6���-���p���sI � IKծ��)�U�a�j�T�{�ek� ��Y�_;t�M�Z�L���i���e3	)]A/�;|��?�P��ى��{2�H����h�n�D�00QK�Lm&w�=��� 2�~N�Z������yMj� ���٢��AX��3�OcY��G��~�F�k6=��k��-E�U1��1�맽�ۀ�ݿ��OSu�A��P����U����IU����s9@y�[X`���۩�`�Iy�x�.���=.�\gu�,u�oo7�7��=H���Q9)��p�jh�XR������)	�(�j��DS�i��:� ���j�㳚��Z�Qů�+���n}{�8顰h�}o�����5�Q��3N�GL.'~=O��*�����@%iFFizfP�>�~ke조�g)�w�7������������r���C�?,��<�:~2f\ic��+fچD��#����m��H69ZQ�Hf���}��5��G���OH#G��g���%�H�U]��SIQn��C&�pg ��D��Y��{-�~�a-��䍞�'!3@N��4 '��%���_�jN�j���D�e�_���Am�z{��LBաm<A�l>��~���w��"*=�v������QU�$2�(��cƟ�u���wg�bT��ӧ�����1�9������ 0I>�����ם���������6������3��ez��G[,����ݛ�x����q�׾(�U�[�ܡg��?M),�*�7���L�q>�c|��N���j��@ ������㒒�'%?�H|VX\�:=�2)���Jm��>��=c�w���G�4Z%�w��'�(���F��6X��M�θE=��3�M�E�ȯ�=���j��e�V�1jpn����8^��a"�Ls`7M��Z�#y��?;�~ÚS��`���*�� ._+�R��PL#�yY���JJ�~�c�����csW}�6:�� �]�*���B�Aw�E?}�o�� �Z_\W��q$�w�B�˹��n�F�Q���a
]�����։�F����WQv�9�HU�������/UT�u�LN��C�9W��%��\5_��TSY��>�/�� `^��5�wSԞ-�_�W�%Ri�vĴK���7��P�=������4�J��zr��c�E�ȇ�_ذ�/,������&D|r����^U����o�t-�-�)Y���u-�w�s[�Aީ�`�㼈Gx��م\�;f�\�3��L������ٷ���?�1��ia��y禕�0��
@�pn����Yl@��&Oyvzr�ZDV�#R��f�*��1�w���j�!r�"W+q(:A���eV@Qk-�[������.�u���$�7m4���_�1݁"�P����y�a�Zdem�7I���n�³)Z��2���4_e
	�sN�m�^�.�CjjCW�nm��+�}�h5��N�j[���凢���	a���ǫ,m���K�� ��IG�y�J c�4^E�T��ӪV{_8/�H�7:�Ǡ�<��᰷�#孩\]y��4jd7f[KI^������=ԡk�g:V������s��R��{�,�D�c�����g4�n�X�k�,B��DI�[1��,h�����D�T�נZ�2%����9��*q�N띌a�
��?��j�nYP�q�h`(3SD�"`�w,,N� QX��{��1A{(��G/m��c�xUPv	MMM����}ʇ�˟J�̎�qJ�e�`w5�p�T)��~�8����[��)��I��h��
��AӮ������[bק_���į7m�d����nN��Ҏ��tƑ�4?��'(���oOÌ����$�i^�V;Zf�>?br�'o��gB�3��'� +�]����K0)+%z황*��*Uc�$�2��i��]�I��,Ѵ#����V��F�����SD`�t5�i���ԡΌ9c�#�7�幖A��QOTtƙ�5NQ�J�9si �ʀy��Th� x9����t�aGQUj�Y���/�:H��� Ĥ|W!4"�TUᥛ��z�e���?�!!�E����30{5W���Si-=n`�ۥ3F�����9QF�{���� �8�NK�>Vk�y����ㇺ0�-ӭ~�bG�$ �:dr�4'� w�m-u����G���4\wg�8����y���>k��x�3�ǃ�@�Ք��q�w�rA��T0~Vt�Qg���6G���(��O�U�����y0!�6�ݧ��e�^�^�2)o~�U��Zм5�4Z����V�����$>:��4V
(��1)� I�H�#L�`��E�Ӈ�ڀ����^�`^aVgU_�OW�*�Jޯ�D�F"��OSo�R�[�Ј�=�v��%|�|��Vh��މ�͖5���¿"o��_$��Q���o�v��!Z7�H��S�/�h�C���G���ju�s<I6;���w�|o?iv���u��T�<m^��_ ,�\�W��f����o��"0�b$g�����6�boP4^+�Zsb�W�^��_� �?�.U��W|n~]ON��?�"&�5��j���<P�����"���K
��,<j��� �(E�aFL����yj�� ��a�C�U�s��x����M���5=3nۈDv�AЖQ��|���K�9�k5��wh!i�z\lu�v:��ȕ��Y?��l,�E��rk��w�1c<�p�T%�@\�&.���J���Ʒ��!=B��^�>=	y��42H_�[���A=���������&�
�Ne�������=��M�.�at�J�+�����q�1�w ��M�� ��y(ߢ�5iJ��М,����p��.�H�	�eC#���	n���,�W����a_8#-,�?\�-�!��U^�o�(��tȄl�������6|�I:�Z�{�b~ާ�-�`���>)CA��~I@�LB��D�������g�d�;v�lK�X���l)b�Ԥ��+`h��A~��$Ŗ����ر>�H E�
��6�8hć��.���0���ݘN�d�Ii�ޥ�cV���U�F�����K�c���E���H�M�m��a�_�}3�۰0(.�C��!�m+��!��X�v����ج�}܈_?�_��$�<���(=w��漟�E�����q�n`N�.-9a��?-�/��Z� ��3����Ɇ�.����駤 �`���U�Ӊ��*Q����%�B��-|"h``�z�h��Ќ	f�x�i�\��ޭ
����ڻ�g�c3��R�L1ݖCKZ��U=.
@�ې�Z�����A��Bb��+|�C���C�KK$
G:��h7�׷x�b0����@�i�nz�v�a[��c��?(��-S �%��(�<! y�$���A�!�����),����] n�~�����?��@V��e����.$���ƨ���Q�3W8`�g����κ�)���`O�Y?T��X KF�`6^˴ ?�v���.&&��+����^��g�ysz�n��Y��E@�2A���2�^��p�>��m*�qNZ�"��k���X�����j�E��5�OYw��U���<��@�M��f�F��Jĕ�5i�f��Cp�-�N!��4Qx%h[��2��V�?@�u�܊�%Qt��_:����=���ZXD���fA\¼���ʀ{�T�T�Ϡ.ֹ�C��}�TQ��ώV専?�=�#�3z�W4��
ű2X����h\��9JkVڡ(�{�Vx�ϊB�Vx�M[�(���x�k�β���e�0��Sk�����y��Yf5���L\�q����Ќ�h����b(���T��
���}�M
��g�+��B5��h8��	�;�q���(��Ո��ۥ{$Vim��3�N7�4	���< �C�!��c����	ߎy��G�OH;Y�3皥�����vwu�� ������8�������ɾ&�ed�<<���Mݴ�@64�"%��+�p�*Q�����6v�g��z���+UcyT�P���z@0��qr������)�P�|�< ����~�a%�l�]�ݟo�:V��D(wu�DK���Q��#�G�D���ߘM�	1Ka:w6��b���٤�VӔ�^K�g�n�0��}�����f3	o R��J�	 :«W^}ά���H�N����b�/raqtŷ�T�\KG'���Kt=�s���>�(�S��h^?��G�5'����@�]�^VU-}��7�~DAf[M�kmںv�g�Ry�����s�IRn�O�a�;"Ǆ���fE��| �@��s���7�&����sQx���� �Q�&�!1������ń�����%�H��Ɩ�}� x���DFY�ҵ�K�
��%��,������ͯ�|Y���\���a~~>��G|�Լ�e`�k%����d^P�*�6!�~���A��n}� ���r���$윙D�3^�n� Y��q�~A+8��#��`9فEXD�1�Pk���p�߰0��k�V;Dn���y�]9_D��x��G[�į�_8�Y@ht�++���s��H�+��yo���k���b2e��.�H���D)9��
��g�����!x��a�-��W! �H;�N�Cn5.�^"g��v�4�A��T�R�lm,�S��ݭo&��s�;��B)+�i1��ouEM�J8�ѿ�c�# �]����p�����cW�����u�"��7%�μ?`2s)�L>�*��=�������R k��ja���� ���{XLLX:}b"����ػʄ����9����ukd6�s�Fgܩ�H����u��/.=w<������������m�H�y�<�wU�OU�>���Xw��B�d����ŽO�*�nҭJ�9[�=����d����O_�'��\O���R���|B���"���=䪄Cn�H�L:�ʈ�v��ѣ�j���B�y�o�(i��Wl���?Y욡���<G����
h�c��Z���I��֦8���@���gzC��u�q j5�Nw�����o��Vhp�O�=�
�D�0�t�hĖo��t'n5A��^�3�)ƙ�Y�[�!����F�oO�tp��@��Y���{����}�^�J��T�s�f��A�w�F>)�
��%ԩx����^�u�����-QWlzKo60x1��\�DL,���ϻ򿳃vӐ�� V�IyWgq[di�e�?�a&zyU��mbJB�)`_i����H�O��tǅ�Һ�w����2ib�X?Xj��!{��U�W�%7�<OG�p�Ϛ�e<qMo &_X^\x��5;��O>b��0����/��m��d��'6�1#'�Y�|!��	��3!�����C�f͎��@���Oޮ��D�{�{! 6+���Kx��o��oh�ZJ6���N���6��~{�L�DV2��)�b�l���tU�����9 ���e���U���.��Pl��'�*���"�'77��V�b���_����m�	��Ժ��!A�l�"���@�7��v�wU��-�?���D�|�	����uğ��f�nB3��Kz���<N��2�f=�i��p	2��B�$��)�б�k�Tp�꟝��ֈ�����s�۫�ܤ�H��,�X�����:���]�����.ܳ��
�����"Z@�9R[^� *f�!ݹYSV�����w�?yb��z�7�wr�Ԑ��>��Gn	=�q���G��o�����>ee���+�M(Ģ�	u�H�_az/�ZG�����2�0}�\�B٧<�!��-��o{���qX�*�h�#_\�q��Rz�3�n7&7���>�+�d�
���;`���W���ߒ��-Y'�|Qػ?�o��_�g�����`M������He]݊����1H<����_bQ��ɒXe�z�:1�^�dg0�V���P��<��}L^T}s��u_�3��Fd����4s:����6JO�v��[OZ1�W&Of�Y[��{���F���~M���m8� � ���f�G�[���ɣ!�aa�nn�Z��jm�1������Cۚx�:͉O�ɛ����G�wj�;���8^�B���b��6��s��f}'�3��b:�(��LU�K>���c�x��)ͻ>wvP*�O�Lh-�~�������P& ��2nFUuJ���ʽ�9�i���ʐ<��Zf6����p��^� ���Y;�h����҈A��l�r���1զ/&i�6��6�?��8Nڠ�}���˩qW�]��J�<H�间{��ɣ��N(|���>���E�ޣ~�?:��;x���o��gk�x��vŌ|��͋.�ة��h��)mFɳ蝯���B����������7^�kK��:S�֪(�2���ܪ�|9���Mi/��?����]tyE��0��2�/e�����M��[_\��{aq������I�z��/�."v�#g�|��\Z��)�+{��ߡ{f��\��q�S��+͉�x��ZS��p����Y7#�r�.���D��� C[^43��_1�ƍ0�����7��iڀ����A�<Ԑ~�r�����ϗ@�AΈF��U�ѩED�z?М0nN. w�{ﮘ��j~��d���s-�*/�H���z�ޡ��ba�_��^��G`K�T-�B����dr)�|�X%d���T��?����3��]V�m�::1팤9����P1��;V
'Q���l7.V��	E뷓0I��Nv�}�sA��ެ3ˣU�O_5N��c�m���[g��=��˷܈��p1�ysr��_��|K��桋(�� ]>{�=������{T���ZE��E�h["�P���wȴ�P�Β>�C|
���5m�=����>5��n�/����Ϊ:�q�m�ʠ��dM.5'�J;�ǧ��y��E�=��_��{��,h�����̢��<i`{R^�.ñ^���f��X\PP��ݡ�]D��Z�V���f��}���v����^56f���.o�mT|t���{m�њR.xqN����}����t(�YV4�,f�C�4���ȇWRUu/M ��| qd��o��cR���icVAL�]�O�8|B�J�6�U�ɲu���\� ����vt��{���_�}>�O�D�G��ʵ��UF���?	���ڡ��-�МwW��D!�������'�1?:�d&��hZ���l&�kw�(�@����=����"ö(�݃��J��9��n	m���G8������S�\�瞙���seu���t�p$O���;m� ��]zܑ�������v�Z��d
�ޭ���-��$�m���0ϏD!�m����	�
_KKˑ}�rO>d�>v�s��٪ sOK^5z97q8Z3�0�"Rg���m�(�x��#�z����	;��_���6�T��Y�t��c��[�&�#�O}�7_RϿ�� ����rƚGI��m]r�m�$K�8���F���N�������"��`�	���cEG��!�5g�l4����O���,D֟(��'\A�Ū��h��,��k,�J&	r�ǎ��� )�&�_��$�\�w�9��t��g���2�˷da1KV�f(�����b�)�姞�#`*���H�e(�����W�>��?�#EG���������5.g]���zR�y���{�G�vV5�7�hX/�s�(�����kH���wke='�<�-�-C�`NH��V���o��O�w�ӌ�7��Q�\.�V�1�KK�k:�!d$� ��F��E�v��[�+r��M/����r���C�{�9�v5������n���%Χ�����L�w�{�����-��l�� �H4�@e��TW.�Y˔�:n>�����t���OٗKBC�Șb���%�t��UU:CCC���Jw�]f8ѪW��η�2'��A��2�Zz^��+�Q�CHB�mY�qѵ�U�f����7#e����i��?����0����V���1��T���OF�77�q�N� #Q�������z4znPlvP���?�z�CAJ�?2�c[8��u^�w�$Eu��������$;�j�:���hek�]��A�F8)��L��&��.f0Y�O�7Lo�1�"W)��-'��+�X��n��7��W��:9��l�v�l�{7����8�ʙ��Znl_ac;������⏒����0�G����,(�	��G,��g=�w1�(�@�`_� �A��wI��������sA��P�H62
���'L>�j��1� F}�Z+��F|���4�9�\��K�3E��O�E��U6�s��yJ6v;�N�~���zl'�����?�EC�	�� T���lI����'��7����O�\:�{�;�� ��g*�Ouv#�	W�,bg+Fh��G�%j��.�~��v�	z=)�}�LN5�g�Dz���y��ӏ6��D�������/.��r&ޙp]t��p�-|JY��q�0~2���,j�m{��n2�,�CM�Q��}�H�oq�od���\�?�����5G�i�8i�+?�:ې8$�8��ԛ��I���j��]&w��0xB"�؝�]&(������{��&]_�p?�S�)K�M�KT3`$�Vf>�[3\ lB������0ޤso;��@�0��:�Lo�Ѩ���c&!�q���|jҋ�S���N}i���Ih�ܳ �T�	*Td����>�6'�Z�V��Z���+Y�/����O�ϢEA�K��"NH@6�ʍ�U��1� ��㩝w1>rM��B�11�?LE�j�Q|�8d�WU�:$��s�	����w�S1��g�3߾��_)K/j�+rv;��,#�K�r�D�Fl��=�9�\d���O8�C��������r� }�uO ߰J����5��c*�P�Ig�j�S�(:��2�����f�O��R0������|red������՘Z�>���MȖ2(�Wߴ�>�x�:Z;lja�{�^�����_���Tp5;H���V��\S���h���I~��/r���r ��y��\��m1<�z��p��!6�|XG��U7WegC o/��D��O�?y<!E~�״gn$�H�? G�������K���EE}�QI�/Z���8����:A-�m�������܃�욒P�Y�ʙ����:appǜW�@O�I3N���B�,���$q�5n���A.m�)�a�gy�U�)I>��ᣟ�CT5H�m|t�j��{ �D�� ������օO����'���I�+�|�ĦDa��j�?^H"f�"��s۱�/�[�J�:G�,lV��T����k�G��ÌH�^*�r���{h���'�^sɞ�Y����4��R���K<s�%��V����$I�O��٧���#��	��%
��؟;?[' lM��Ӧ?)��x[[3�	�Q�u#i:Nwj��]Cic(��a��$*���R��v����A*h�Z�&H�o�$��X5��
��_k�6��`b �I��q����3��؈�{Dܗ����E���=65���)Ȍ����*VY�՜�F2SS�����ݸYU�щ)�>��*��������U~;A�����x��������IV�Q	��U�~�OD�v�$��,V�3>A��KU 3k��d�9��k\�V�Ygxۀ�!����0v�
��� �q���r�OC�.@�� 	���$$)��َVkݮ��]2h��֋�<���E��0�#{4e�:���gᰟ�B��b�V���SƽtIK=���p���M��m�����o���r��a�M��	��Ah�x�Vt���U�͸��z3�,�B=��LE^}�h���^F�iq0� �}��"��0���Ji7���v�H�R���G���׌��F�/,��-3�'`�*s�U��Տ�u*>���)!e��`]��#��d�$����!�F;)}�H	`�!d�*x̠����^��	�ʲ"X����i�jR��/�x�r�����F����=������l�x�A�<uӕ���#MӮ�s�UG���� u��%/(���I��6��T�ͣ��)FF�у��c~z�X=A�>p?�����K�1vg^���N|��]�@�)Ƃ�hl w�R�{���
<���0�y��ۍ����&��n�<�����f����3\؏�����mVe?�n�#,���ī��^�pخ��,^-P���e�oW	��.*�|���T�� ؖ��t�o� 0pb�����3B�2�W!Ig�HC�����D���' ����8�7g�}f]��n�%]��{�"�@�q��� ��7��u�8�Zj������FJ�'ϢY1��*C�n�����nK��Huτ���;y��=�MOѡb����h������}]PR.x����&�GD�\u��d��P?r�Z?��7��;y�4YY��RX���K�BpbŖ��v},=���n��$-�w�A�֧����رM�-t���i"������Ǘ����n��G�)+.�p�������{?����ɵ@W`��\Z{B�{�q1��<��������`���<� R� �V�Q?Bʨm���$���=���ksH�ݬ�����Y�(�Q@�u�Ƈj��{-�tH�Ů��`̈́�E�sJ���ᴹ����h�sJ�;���ww�`W�u�]�X<�'E�r�������0�����{�pa�4�يk�O�X��!����n�PJL
����!�9Gp?1b�[/�v�G�w�n��OF�"8��e#���r�X��7���3��l�a���>�����s�AwRr��t��q??��}.�\i��ܛG8D�}��?�C�j�n���Ir�3��m�����귋�+�f��*]�D w"1d$����U�'p?��P��j�Jg�α�5��H��c��x=���"�ݞ�08�^;�p����v�}E�Z�Jt�K�V/�ra�3�s�@<�A�1�����[�%K���2�@.s%�+Պq���,$/���i�}�ȞE�?5~f!�^sa�׈�I��2�G���� IS�FW0W|1���_��NHM����6�`����)���o�����'YD����\���x�>��T��T�D��=+ۑ�i)9��^ٺ��D�p^c���e�Z�� ��9�KBl���b��l���zf��{��'@����o�}1s���a������s�:bu�<.��MB!�M��!3 �lz������"rb���Бs��ˮ�l�j�&P��_7HKNwIJ&]Zæ6�����_��L��gU��*��3�d�f�Ւ,�����W��+�.�g�	���ql'��4�����RX�3�.�z`�~�A4xk��{;�%� �{�����vB������V�{�g|j�.�����
�w+��9B��OE��/���V��!�_T�q�b�?��>#�ȉ9Yy��A_��͖�EK�Y���L�l�#H^�<I'2�Qt+=���򺺈�b�]�(GEy&0��z�ex����k�.�*`4�j��3�'�c���>����h�:(8%g$9g*�F�,�s��-����{�l�m)m"��x��M�9*5(�r�T1X�����S�{��0��8����D������g�ȭ:��� x��e��Z��0���@��>][�wh����ȴL���ؔ�c�G�	l�$�pTOD]WOk��Q�5�{�=�R�*n_/�6X�V}��"�����}��x�<�s7���_O�bg��E��+��$��	���k(TP��^%�Y�T��P�����y����e�oא;;e���(Z����~���
�8=Ӯz��P%�����Ɖ���!����N޿~Rb�<{�`j�?�k�.%b��f�����2V���7��O��"�p9��EkOo�:El��pN{�d_���G�.�'���rk�4�a�9�+�����Kb}�n���DÚ�:�C��"}��DȪ��S��O���o���>�쯥9@��ٶ�ހ������Zu��$!�m5/�ϐ��O20;���iɾ{ܣ$����G��lv�GrGeUy�6�J�P=�q�r������Hv7�<|J����n^��R��	1��K�ĖR��f�5��Y�=�e��'�x�E	��{ɷb+�o��H��I�TY����.����߈�\J���Y�b!��ҀOt4�����M́�s�ǹ��dw�r{����"�I�iչ����;>+�z��+8��eH�|�Qא�6<ᢑ�asx�����N�NuO�~�"_������)�ҧXL&��W�m&����	ϋ&5�Oq�C��j���.�w1�-��/=qX��}���6����~��e��ߟcW����' �n�sE� ���}�o?�o?�4z=�B.,��ƣ�Ӽ8c*��?-�?�B�����!F�xD{R�(EHZ8	��1�c�lz��{P�O�4�#������4���}x��т��?�s����Z�8�c�So���r/�0�wXW�Q�T��Ru��*i8n���{40Rk�x��_�*��U��_�]�K�:����LP��e�3��m2sɮ�:>
��S���8�H����͐�]#�`R@� �C���=�v��^��~��R
�>�������^
2�1�jv��Y���4�:?�XE+�/���`ȃ�מ(�����>�A�_ >9����z&$���>�%	��n:J��8dP������=��'��S]8띛{������oG8��- �D�4h����N��E�5��7��Ѝ�o��!ϙ��)�`���ڪ6�A��*��1/]�/	�
�~[�K|����N�$q�*XbG���4��C{5�)*��R�E~�W/��I��'�<� ٞ���0	ջ�m�����5P��Sg�)�Z%����o�:,�5%1�7X��9�q����/x�!��r��sw>�5� �@� ���z�Bdf R�[-A����X��ׁS0��%:�rg%]�����9���-��U������ "��Fq㈏�ذ\Ҩ��<bټ��sy= �3bI�pU���C�*]xy>�A]����?��w�15�P^��fWK��/ަ%�`tE��!r�Ԅ%?s|�t�H7�h�11�=,�H�� [m����/����L`T�"��uK����/��>�KZ.9E��Y���2�i�u��}��D�:�v�w�=2� u�p���E�\��PXY�w��}�x���v#��<�-����6~8��!��H` �EYJ��,�$�Q

��/�l�P��
)棨��<��$n��Cey1=�ZLX��V��ˇ��8�jNe}6�b�� �uO,���r'� �8�D�~�)���xT77������x�A	���t�e��4q��x�Z\��<pt���z�\�i�:���������k�#�o�U%�GN��K�7B\/��
`��?����=�8�h^O��?҄Q�9z=F�"#�g�Q���������z�x(���V��$�t�5��)��-�9H��4*5�Ց������SMm�Q-������X���z]w����������~]���z]���tZ.�M0��g�۫�� ����E"����Т�AġFպ�u��6��{��sH�]��F����+��p��L�<:r~m~>������䤢}�¬�����7#��;�e<V�>��hD���:�	r#���8Ht'�$��x��!�t������o�ʕOJH\��mE3�{{S&�ƍ��L�]҈�d����-hq�t��^��{�_�-7?,,�g�]�4$�VP(IwQS�[�+�>�]�k�nb)}���/~.&]�K& �/�l�f�~�r#c�^���@>Xr��it����g�4�3\��M'�xH��P����l�����_�1^~w����*�mF+{��\�@N.b���]5v����V@9�M����#
9�GR$����fD���a��4Ĝ��Gg�?��x�c^4r��%��@A&��a�i᠄�X]�88	�p�Lc�<Q��b	pi
��U�oe��������{y�OJw]D�C fk��zm�Z�>����A�]��}��g�:A1w��Ee����^6B��I�����8���ؿ*YZ����`����E�0Jg��L���J�'0-��ʭ
�-�n-����Ȭq�ԟm7k�cN��u�$�KQ�
W�j��|(+��*�nLw������cb���q��Qp
�3ޮ�Mӎ�ɩ��Fc����������`�S~w���m<~G�n0��,�B!/���ȔLː{\��Dt�q_�%���T7^�<�:Er�	v4����l�	eq~�ʇ�����K�D�,y�,�+[�"��YO�V>�|5�\��x���N�� Ρ�y��{�v�7�i���Ga���ܵVJ�/2��F��W��u�����&�� 
�9�����B}@J�G����!���O��Oz[�/�{���9��s��X��B#�p$�*�v�x�A(
�w֧9��I�������ޮ�Z�,H���<��]y�U!���_�ap�{��b�=�B��֞��a�aM�Z~��i��O����r��6R���E+��K/L�xkoQ{V�a�%b�k3���C���9��|�i�ŝ��Y�hX����N��W>�J���V�t���U���YQ��l��QW��vZx�˹����j�Q��D��)���6����S���vn���Lqbr��������k?��Me@��'Nm�'����R?�v}�_a�W�d��[n���:���	'=���=������U��^g��8�bU�8A�(�ȿ�0��.�WK�ޠWz�_\��v��>�YW�X"�Ѩ������L~�"�J��p-��)�d�"�!{Xc:\?s��yÐa����ǧ�6*>�5����qS-h�ڒ�B�,FW�e��������wc#.0>�<��o�W`jl,^{���%QkM?��vK�!?��H{�q����Tj�p�D�ݎ�{�M��2>��x۞f���&�ˎ����ՅNx�ۚD���$�d��IF��×|���q�R�T�Fc�{�D@cЁ��6�\�6VG��Y���q{VG�z��	s�c��h\E��r����v=�a������b?/�<t�]��-�$���g��POʝ1�ud��u\���+JGV!ҌG�O�����+��ri��z�A���&È�\he(J����Q�h8����1ΏͶ�8����W��6�!�֤�����E����im�UL��}�1Y�N�pk�~�d�ڔ�Oca3��Uh��o}��*&�ܴ��'r�Q�i{�|�ܨ���0 �G�qѕ�c���{C�Y�t���!&�Z"^k�
=�k�f����*F~*�&e3�8��D�y�d?���o��re�K���EeM;G�����,��Z�o���P�c�#h&	#�R~w4�OA� �\d��)��|ъ��+J���/uE��W�V�j�3j|I� �ױ�TL�t�i�����6��Lh��V7H�^���D�z�#a~�8O��RO�
��⅏k��],P$׭(��*ĸ�v�_Ǟe=sƑ'�\�S�>8��W�64���&�f�~�o���x�6`����~aW����o�	�r��"��p06�b��΁<6��N���Z�?�x�H ���籓tؽ�O�Kw��Vso��둗�Ak��3T�rL=h$��)����nN���m��w�����j7|�+�O��A�B���~zg�/����dJ�����BaK ��8����ӥ��	$�[_"LD��E�W!��ςcf��D�`-�i�UL���]OD���Y���9��m���\P����X�L������*�����=~�̙iCF�4�I��f���Z������:���G����Ao��U�ϫ�GMe�n"C�V7��G�_�
��PD��ƒ\�g
�pC�RqX
ڟ�hz�,��C;X8��y^��\��D��,)'YC[�Iw�����ze���S��[n政��u)��<TL?_,���2J!�z�y�� ���Ӗ.Ϻ�,�3��d�	�B��r]+.[�л/�mCB�������<���r|�L>���/��],����`=M_�.��ր������^?��ڹ�` �^2�>h&���q���P�x��g�T|�)vy>)��6$EUwU?�<8r��Ϲ��uف�����^�MYub��)Po��﷙N�o�AK����@��Ӫ�(���.l����%�/��,d���Ki��*�ǣ˙\��'�L2fY���*rҙ���T2�r���Q�t��M%5�+��H]P�Dk�'�ݽ�vJ��>���U'*WP�.����/�'�DL�Mj��)�z���w�]�d�0�X���Mqa`e�ߵ,6��w��MJ�����c����F��YW�S��E�?=��3����麌�Bk=�K�.+���wwe�UOπ�@�?��`M��Fv�4C�����^���o�����e�����6��%m)�E���d��⒔f��}L�ɍ���%	��UM�ؐ��y�y3�@ꒁoI�④r�UZ"��lAhr˔�x�]q@yD.h�@r����Яx�t�X��͏��������LL��N[W*����\he>������0�yd �!q*/9p�o`�����*ab�bBr�?V4Ϝ�M����37fZT�4̦�Ӄ�L��g�]�9��o@��)��zZ���\��R����w�y�h����v$A�x��<M%A���H�H_Wi�#<�z�n�Z��>�^ɸ�!X�'���o�jW�~}r���m��P�4-˛.͏`3��+��L��.]I��q�F��O�uІ˞]~�L�W�H�G�.&�g���Zr�zzeF�Q���ۄn�C���*�2?�<��g�Í����H�%)(�-�C�1�#��E�e8Vzd�^l�5lNo�G�J�26�h4���I԰E�
�lR�xq�Ir�^�Dnr������n�{5g/����SGn4�ZŽo[�_v÷.=8e�c��nu6�"��X���uA�A��"��f��EZze����~4yD#SoBn��wŝ#[��#�*��y�%��Hr�.A���f�\����W-Oו�`���@�9�5)@������(����~h���x�?�9<���'~�!���X�W��M��=Q~�*�=	�(�}�;)=�Y0Q!�?����~W��p�{ދ%�ֳgh�D�C�T9{��nF��Y�fZ��N�fǪX<���2��YC�=��Q̺��r�N���8�t��G�Ȫ,;�[��8�!;�QC���UO\Od�!�n��cAt5�7,���Rӂ��ZW_|�󯤴;��,l"�XiT�͝�Q��J�獮��Ωx��R�М�0"�{�F{�TŒ��qV;Y���hh��vs� ��q��N��E֔��3s�j�6��vz �٦H^�$ǆH�����W�>�X��$�����o!�W�wpQ����ug��K�ckrq��'�����zyO[��?L��r<9���7D;^�t=�5��n���d���lJ��OvͶE,���I�v�&2���U%LJK$-��I��������U��*l�/����篏k:"n ׿H�]�o�\��~e9�M�%hA
�攔��з�i�뷓b��A�qg��u	��awY���('ϔ��v�]�4��/�^C5��Yc=�ˍ��U�U��DC�5)-��B�**ý�h���O1�'�{�!c9��������,�c�)��yO@�Z�&���0�2����.�J4������NCi����Y� �-�^v��,�IvM�ӕ�c�ߐ�)�E�v�ʼ���2�'���Kʎ=�D�P6�mZ_&Z/LcK��6���vM���ZN��.�6ym��\��BV������o�}����;�ci�Ip��Y�n���+,�l��|	�z(��r��|&+������q�w�9�G>֖uس�̠�Y�)�ld��rM��Ӣ|��_��K�ݭ	#g�~�`��N�{��]������]-���{?��К�tK@�6�h�K�9O��U㲗SEO�y+!����z	J��q�R�h���O^C�d��&����c�5��M�?i�r��9�|�5?/�z6?��'�\פ(�ޏ���=�Z4�hqLJӌ;��#�Wu|<W��Co���`u!LpSy�y((u%~ԕ��Y)����" ���eM���r[\�3�B�2b��K�`��t[��`����.5����f����np�+һPD��ۧ�i+K�O�aI����!T�l�,M� h�fC�4_�S��4zWS��N�_C&a�G.o��߼$_��VwS�%��4",���0�c�LB����X�zl^Ŀ})��[�50I[���\�P���~����P&%®V|�)����;�.���;�X6Ò�n��=�����,�4n�U�O@��K�ܸf��C�h�/ٌE,�Q~l��2%��cG@����������x?�A�A�X����2��A��Wӟ����Cs�"?}���~�������H���D!��~�b���%��!u�h¬���؊�d�6�QG�v8��{��;r�d�巑��������썻�OKN^��B-���vUBv6�n���e[FD�eee��p�W���iM[aQ�-_�eQ�W�|Jb\YS���,e�?��.D��422�#��vy�$����k��^�2epy�(YƗ��-�%��\CB&�\��%�mc�;h��4�#��`2��1%���(�Df!��4tM�Y�ocW�n���|}+�U=zT��QP8����N��%,�Ϟ>�P�=Z�����ۗ��p[p���XDpx�Xz~�����΁-��>)��VU�[Uz��I:�~�GȻ�nO[1��M"c|@�"�R��疖��4vD�@�#ig����v�c�����a�E8��S'剸!�GC��MU�ZS�eK*5Ǻ�t�%��d�"0�0��3���*پ�.>]������iHK�Ӌ����u�T��!�k�!Q�j�=E��N2j�P.� 9����@�e��V�p�BL�ړ��

̚t m?�m����1Š��}>���6�.)��ǓǮ��k�y����K�R����D����0�ӛږߙښߙ[�%;VP�����7:���%���w��lVRh�ҹ��2�:qִfgZ�RYO6b�4��+���Xa[y�g��zDO׶��b���j�zudb�^("٢�����\U�;$�c�����y+�ZU���&zjs='|�𱫰K����
����;[���b�+'�������q������	Y���b�	M��??;���k����m=�+ѓ/��*�n���;n<���_�ӦD)..{��c1J��CI_P�Eq>�ۤg$]Z��l�zX�J뒉(A�7w�{Tc(����5&CH�6�m;��P.�#W�M5���/3KG��|�e�a4-���1�P�rZ��K�!���a�����'��"/@��Fr��;*e=�R%�����Ȫ�)J�sl�.�)�ƾ��h8]����k _r��8��yJӗ��W1���q�vR�Ga�5j����Au[I�yפw�q#���`�t:籆|��$�IŻ��|���sy��'���JK�:KL���ƙ��P%a��*H�=�4-�D�DJ�����ճa���5� ��5�Im�G��
�lQY�W�|Ϭ�i]����G���h<*�7����{4ȫ�,��[l��}7�0x������Y��4ׯ��p:��+~�pě��:Фc`�Ԡ�iP�������[�����z���f3~o;�V�$8Mao,��iA�D�ܦ6��Є���e4�ee�I_�%޽�pz?�磻�����K˫��m:�4���'-{)�!���1�H7Aط�R�0�LB�y�f�z7ɗ�rz�a�,$�����Y��=p�Mv��m��[58V�r9�N/_�h�ݸ�~Z�L���4ޓ/q4t����+����e��@�\�C�H>��t�w�AOJ�@� ���X�p|k���ɠ��jd���(J7��l�J.�u�y��	��F�X�� �%��ޞ��U��&O#DKx����V�m���:�O��
iق��,�mC�f�C]J�R	~��QoX�pB~l�$nxVx��Z�)ظ���j�1��c�E�-/���3L�t��q��=��j�������&RH�8�h �}�ʇZ����B5)���:#�/He��dG�&����*�H�X���g�($G���@��E��x�{u�U��8z�{�m�^�����p ������i_ٛ����A>uho�+��I�f��H�c�\Z�m/��%���c�@��~Cȋ̮Pp2�;k�����?x���8��c���
ߞ�ᆓ2ߺ��`����z3�/���+�2D?�����(.����7�=���Y�����^�L���m̶����k�z��_�,�{��g�*��9�X���Uk��޴���x+��D�l<9KJ���Ƽ� �2N^�X����՛���3���DZ)qg 棭�~��d�~V��ƻ��^�R��m�S'�Χd%�U��8�
O8V�NIk8�5]���s���W��\ݖ�I��(ga�
g�v�S<	�ϡ�\�YPꭩ�=�dΠ���r�3���+�m�P����TIҲt!����d��Ҥ�ƠKܳaY ��ǆ�ϑj�:�B�+|��]�ʲ/�F~�BW�	8�1{/-5����j�2]��`?��яyZ*�.�ń2,�_h\���������D�����[N)�lȮ��,���D�@R���ld��i'7���*�W���>��\���à�$u�	�y�#L֦��.�
��`C�L�y�\� c���ͥ�P�W?�FC>���C�"=�J�ٓ�s&�{���(�WR8#�h��O�aj�$��E�K�����`����U��y�a���涁>��8b6�n����0��fI}=��!][����VR��K`�{/ �G0����z���R?��DPg>���*���O�G8*�;��7XɠkWj����0��$s���?�[[�Υ��K�=Bw ��:����G��	�ߋn��J��(m��F���(Ě��l���.Ĥ�{��qM��nx�}$<�7m]����l��D�d<n�oT)_iڂB�cʡ>%�_0��,*���\HVZ�:�'u&��dL���2�������/k�/�p�dT�lJAQW��e��Ӟ����ot��6_��C�j`+|�P�U����C0p��,"�0����ND�P7;���Ko�7�qM:�㟽��y��fa��Jī#JQ��P�]M>b@>���S��xiR��}�t��,A����0#5�՜V�&[r��C޿׸%5��5o��� ���O��f�=��/�8�w��ۍ�Y��ġ,�
1��?�I��x� Q��&)����Ē�L�f�JE^�Fn2��l����i&��E�&?�g)����O�ڥ�|J��o�-�o��gV'Y�5�D��U������~�խP�\��t�X�.O(�G�%��u_�u��ڊ��y:���?S��{��a��Z3ra�ݍ�M��I+���8�K��˰�������� em�S�.�L�&�����,h�M ���޳�/��^���a��Ʉ;��"��[Nz^j����b/���������Di��>A�YDc�y�f��*WCSX�ZI��ɟc���5y:K������;��S�-�n6xe�	����<�%���7}�YL*��>��X�^�P�@�6�8$��t�*�D��CM������ c�HD���k2!�+)m�JW?͖����w��lM����\!�j5��=�RpI������r4��b�%���o�Fn��tZ m�5p��!��x5�e�Gd߹�E)`����=^Vm�B��pz+��5�3��Z� ��ca��O/ 09�;���I��ތ�O��z�&�W�Zq6%C�oGw��:��2YGpV֌k��F
��U�f�AM���m�(���?�^(�|z�W:�t����s�s���E.����7�#֖O�}P�wd�^Y�����,./11% ��Xv�I8���y�߷�"u��`ܘٯg���i��AI_=`�s�
&�&%6�H8�����ᑗf�V<��OOΈ�"����\Me��2�5�q�Z?�J:^�t�H���A �^�+(`��м�G(�&[���/?�ɊLj� Mbƽ�~4�mN��zs�@E8��5������66֫����_�5����( {�G��p�˕�U�U���ǡ��{77-#��u�\�r�������1	����=�~	�|:�k��PRUEg�,���|��g�^gc��Uw0�nt���:.[\��
����bCy�sZ#�\�>�^�i�!�:5A幮)��J������T��������ʲy�=�OĜ���z�"<ח3��r�JMgg1�6\v���pw%Т�=��U��S(VMn�����t��I�wњ6����1���I��Q٪�����~�^�n�Z#�jX�GD{����K��=�hO[�Yxs`�g���:����+��s�9z�	��.Ƕ"Rt%�{�C���J0��M;tEZ���P�A��թb����|e[P��ʠE(b]�i��\ýϻ���y�F�#^'g�QtT6�T��.׏+26 a{=�,ǒ�5���v�ᅵJ̺�Z�|Ü)DB��#
X�ӽ"t%��[j�#�m�G�G��q��5+O������F�:�{&`o����/�C;���Dd
::��R�A�ׯk�(Ĉ�#{��U~k�A>��T��Pdvapo�����
���x�������w���%��7���_|�����ƃ��Ë����3�L�������b5�fQWd��⡖�ɑ��//Gn�F�����_E����ª�/ő�>QڍF��"��ǯ_[,2�rUJC�/u�ӭR��ѭԼX�5��gC]ݨ���l��fm�fGz錖��ƻ^��
7�jkkg�ߡ��k�ϝ��Q�����_^lol���#����6Rh0�m�-�f��-���
1[�"#��S�;i+����9���胦��kH��x�!�-+�X�)~4|����mDͼ�(�<�-�x�J�PoA}������B��~�ʘ�ƈ�)�IvȬ��
�����Mm�I�o���E~
���?!Y��u��k�x��'��ʘ�O�b�7ҽ�j���B��i�
�٨~�IJ�VJGtכ1���EC>��� p��?�q�_��R�2�6����As�x&+d�Ӹ��W D�����k~R�뢤���2�Q�g�����'��XI��t�xv��Hjg~g�bL�a^m��T����:���������H�ېV�v��8Ո�=ţ��jE��X	81mܜ��5��]Q!�$U_I��כ��'Ȝ,�s���zZӸ��Mm�TV�[ٖ5��i�.Y�Ⲟ�∱C:�=���.���;�SD�(�j|��xz�Wh(��Z"��w��>���~��ŝcf���#V�^�h�d��qz�kZ�.����1$o����5ɱCqI����#y�L��#-w2�?��B���՚��/�^������gq���R�K��
T���t�N�z님&Oqz�ŀm(
�!�D7�C>���{�稙�����E�4A`�\�+�u����h�{&f"N~E�54��ڂ��V�ϟ@�"p�Ho(ώ��ZC^�w,�ı��^�_M��D]�^m�e=&(�b����T���q\�'4���Y�Q�ʥE/�m
����+�A@\�>��U�`��]`12�u7���y�y���/�����%Ɗ|�V�}�V���/?�Y���T�k%��`X^�U�n���v
�=��Fವ�t���w5W����D�qC]��
JY�t�Z�;�;	g��[����B
��m�?/(��K^B.���6��)��c��%�ؗ��k}mV�G�L_`�s9fL�MNcCʨ��ID�#\c���z��������6�?���,4~Z���T�,����1R�d�u�Lm�V��)���_Ojץt.T^|Z�z�W���]GQ���I��@e���gb�3�����`ڳ�]^�?o���g��,��>���'c�5� ���&P|��#��&ٛ3��Y��4�)��>����R��Y�2�#c�3Zv�S�
wӴ,�����ia��R�'�� ��5RL�5����'$(�79�c	e�1�G�Z�;jW����:T1YR�u:^S��xq�P�{,�q���Xeޟh���oG/�Vr`3�GZs	�獮9Bs7�u��\7^?��V=#0��.�R8ЇQ�xP��r��AXM��9졷R��� �\��(�C,�����E��=_q鷩ě=����ej�D�2���{oA{�-|o�}��=�|�s�_�X:��*����C1qu�[k)R�v���Hw�3����;)0�q�<��hM��K��
�5&�Ä�|��uwF��A�a	L�B�# ��Ɋ�Β[�ү��!��E�$D���� sw�w�dH.3d��x9�Yw�7�n���QY�Z�9m��= �������{�uJ�i.����e�03���)نP�� �R��|��8�H���	�iy�{�O<��0T���r�:+>��g�9��~VO�#���j2t�3�2Y�����@��Ѝ�`,Q(��d3J�v�!�L�RmTl,�bݕ�N������w��5�K��ẒR���/�إ�G�h��q�S*�H�����'X#���U>��e��0�#�"�E���}"j�G�ǅ"&���=��{�\d��l{��tZr�i�N�c�����9R(�F��m@
�L��8%j]�6RT�����|�<�莰�'��sD��\�*���{�fۻ��4������];�p��Ή�KL����x������ќݗP��t	�s��X��T�Nƭ#�hsO�^2zQ��rBf���g�6G�F��|
Lf�_����|h��ۼً��"�<������>�F�ai�|޳���i؅��8!4�2�Y�(;��y9�����ĬV���c[gC�O��uF��xG��A[�`��{|zo�L�,��h(�?�a������C��Q(\�zn_�k_؅����50�h�m�
�:F&��5_V1U����V� ���g:[�v�"�����FiYR+�{�J�~��j*a{�i���\��@X<��|̲���l��k��d�������f3P��.����%�5T���#�Ͱx�����1~�5��X��{e�_�����~Y���7�u�l� S�f�ف��8�n�CC��3��Q3�AS��5���X<�G�(5����2�]1��r �X�A?s��/���!�(O����7���]/ =�Ȩ3 �g@���&Ê/�P.�@����L'ܟq���9ձBu;�K"�����w���^�s�<U)��z�l�r��R���[������O��#�{�]�&�^V�Ǆ�����/z.��������.�I��=�+���R�+\oc�O|�3䏝�������_��Q��u{h�J`�{U�����x��rv� �տ��2?����M܋�0Z���u�y�9�����ٝ�48w-1��P!�M�?>�?�h*QsW�X.����x׳zm�`f�
g��xc]w�W��;4��uF��P��l���F���H�;0�u�R���K�*Z�8�P_�2p7����?z!k��a/��|����/�*���I[1��x�e�l&������Φ���|�<ͺ��B��5��Ƴ�E��������m$�ۗ��Q�����G�$�d���r�� ��S����נ�,8���^�IAe�eA%�Pn��maJ�<�Ƥ!��>��Jx9�ķO�L,mX�h��q����wX���=G��T�&*.h�[g���r%vR�pK���K�N^a@L��ݹx%qa���Ǧ��^�^�7rD�/ôgy����Y��NZE���I| k3C���z$:w�b�9B�-�'��l��?��d������7��~g���|i1��T�ҵA���{!o�Ǽ3���m9��Åwm����^��*��'"a���px��k���7_�-�3��a��ƫë��)��.M<�7�z6}�11����Dp[��W��aM�#�+�J�NH@N�%�&�
)=�/�Bܯ��.�r8����;�J�/�9�c����I�⿊[������[|���Y�S�<����J������A4���k=ü�O����jG�s�y�N����>��'��#PrQ��l"�pHd�2^���2T�9���{.�0��K�X��b���,^�����6�J?ieU�U�+��)�� �v_k
Ѹ���T�*��jn��C�M��g��wT�[1�IƄ�PЇYh�tMR�Wz����n�~]��,�������$aK/9�Qfsh�P�$'5�Zjs���I�����l
��<K=j�"�I��j��^4�^N�'�IK�fͥ�m^���lQ8~�]����K3�<ӧ��/Z���ܲ��0��c��
�	:�ZW�M���{�$���zmcf[|����Gr$��<)����Orz�9�|��vwَ��stZ�~E��wt �0�!%���hAi�^a���4b��O�h����m����4n�hY��W��&Oپ)T*����kX��[?d�S�����J������UdDٹ���p_�"��[�W�1�+��%��-	.*�ώ����A���0�P���n��D߫������Z�#�����GF�7<Ț�l9�'pP�t%ɜ�7��lə�����V��A�F4U#i�6`, ����]!��g�rw�B�&��^#ZGL����j�_���ׯ�f�/���f΄?�9�<>��0�5�P�ey�)"���#��#�#�m��_{����4�@��љ�Waˊ�d�Ee�pgA׸-��]�2�����N�!�7ލ7᜔�Z=�7	�nM]ITӴ,*'Be��%*���<zY��YH���_��d�P�JM,7��30"�"���"�Zq�ߠ���1XP6�_=q�zҷP`j�M���c���(��r��ğ��ii.�U���_�0�����%{�c�j������"YgA�渦�l�=���x*!6��6��1��þJ��&��!���ٰ�{4�/�������N|���$�xu.�k㛈1�Ä�5i��R����~�<^^�Ug����H�\c����9��i�U�Ec4n���i��
�41��� ����!����TY��B�׳����K����)��!��w��T�5.�)$��d����1�S6q�7Ux?�m�<]��?��,�plp�j����5����%�.ׯkKhcT�s]�	Ǉ�R�NfJ���( �6�G��5�G��U���E��ض-WQ��mꆣ�%|�H�����?�X�����#U������A���-*(�56DN�.�H�7M'����'����x ��W�C���ׯ����D��
�$���S��`I�f@=leW��7l��0�j\�|c��s�_i\�~E��M����OL��������� �©�}ʞ��H�?��u.İNP���M�n�R_�r~�7|�zŉ SxE?�蔥T�t�eZ�y$W�����>G$�J"[�(Bx'>V3JR.�C]j�;v��&����NzpJ�4H+���<n����A�Vh��4R�\�'��^o$ ��gr�ޛZ?� �[��$�l�@�)��/���s9U�$���w�뾆�[#
*�.�z���d��t�4������*�g�@$gnῒ_�g[����P�\F�f�'�fD�`J����uM��	��v��1�;<�nb�Ƈyd6o/�+Ҩ�7��.�c^.ڰ��1�h�M�py�� ��4LNk5�a��[$ܦ��P�o�a�>���Y�+���L �����&����|�3�Ug����Mp�D�Z��N�l�e��V�>��\�W\�����a����9)6�RXDy�ti{����� ���X���L8·1��~4~�:�����Ƿ����A[c�!�]A^��5y^�����f2��c8fŴ7Fy�ba�N�=��	�j�#����[�����{�T،t��32?;n�Z+�r���Z��%�A�!W� I�}�W�+9kg{�^��T����o,
K�xH�ӞaupI�cE��xS�q�mU��y��F��/	u����5�rM��5���A?/���֣8>�eʑ�P]�Z��%��#����Jw!ĸu�����5�����jROƪ��]���	�\&~ GZ����[B%A��g��a�H�J!�������U K�������E3��M��@4�����v>�K��ohÜĺ`��j�'��c�B�E�w5�1��	�7����n�i�a#v�/䰺�݀��W�a\�N=��.`�V�U�LJ�E�ͥ���m%[��g ��xU�=�U.�ʟ�?�݂�w�e��I�Y��� �`�t�9$�A�¹l���PsP:�+����'�Z��5�t�Y?7g��d�|��g&ǯ���� �?��%�=N�bC8�}H�Y�{p����$`��#I8�	��0	'����{1	����l a��iL�,���4 a���O���}�w:��1	�tW;`���>h���i�.*���o�e/MK8-"�4
@���=|����o�g��M�UAEs���tq��g�Z�
����x�ʅp|K\�L�»���&������R���Xp�f���,|���Y��h��<������x:�~�]a���#�V�� �����S�flϿ�f����&̥���Գ-F��b	�?3�����(�%㔰�}�U�<�n��G2e�~�ٵ�εm�!(x�һ�N��$,o,J�}S��=���S���|�����y�F��RCa��X�14r�f���5��*h�-���8��� �з��a���:��/<���?��OK�OS��$��Z{+A���7��(ȯ����v� �}�!;���ˢdP}��%�|�4hY�b�Q�O���)��2%غ��%c#Z!2b?����:�뚽�Q<_]�A+�G6.윶'z���t���ސ0�Ϭ�4s]�"p�t^�w��=����١�|�c{�[�omڒ���ၡI�2���'�ٍ_�H��G����ҝ���_P
Rӷ�sD^4���}dl�l�#�����8I���Q�矐�t�}��<��+�S�?w��B}P��w�d�x_sP>�>o��9�qכ��Π�XJ7X>��>]}�O�N[_q�x;�uG/�Z�k�d��x����M)i{n��wm.\NU�S�����(��)�(a�?.��l�z�o�ɾ99��<p�իz�P��P�z��Ñ�}�P��4fdLqjzB�̠k|��H�SjwQ�t1v)��1Fk�L���?|z�5�j�aC��+��
X�l6<y���C�K�\���;�G�B���캿@��um�\p�{fS�:Z-%W't�/�����S�"UI��$,�F��N�l[I���![Q���Q���Kn������Q��Ypx�F#Рʹ�!�����<r}u:�_��&�/?P@��rgc/"��������0VSK ���<��z�F�/��c��B͵����O�A�:��9 n�����b���s	��va�~h #���m��3���8��&6f�\�I��M���Io���v|��ኊ��q�v�M��� ���L�� �x��~	�c�n����П�#m�͐%����{�c,R7N��{`��p�:)1�d�v���,mp߁'��	�;� HbE">I2��`{:N������4��l�ף��-!:Q�쳓����T��2�5k8u�����j	�3��7t]&�Ґ��B�o[X����xqU�!�3��M�|��OXd)�~E{c�s���e����Y@��-� 
>�!�Ĕ�oJ別^i3j&��x�"(d'`\(�R��}��l`��7�x�? @���<��4B��<�j1
.��!�Lt�y<?;�%����W�zr��e��5�w��W�~�p6�IGR]�.q���*Չ�%��Fy#௒$�Ulۈj��7�����?��ULka)$�VB߫�?�=$�JN�c�803t>%�7���L|��i�I�͡� ����d�,�o@}8�A��� �u��.�Ô�5�i�5\_���_䡊!_�q��| �ngL���	ݾ���͠x�%���6}�f�m���G �����Ed��B�_�m4�Y�L`�{������A�HmȌ������Kg��1�2�����,��;����`C�c(>��
f�C�t��-�F��Sא[`[T�
����� ik�PT��F���̣���s�b+qf��'�������|Cv��M"�y!8d-�����#�gC�U������_ �}u-@�%5�A�����I/Ĕ�C�|9��Sߝ�c"~��qo%[��a|���Q4�o��F�+ޜvZ@���:�WVa����6�GU�l���.ᵱ1���,,/�S���?j����	�b��Z�!�T��e~��0��R	�GwNb'��r���*�I�0��M5���VQIik]��-D���p��ڎ	�!Im�~��ʝ�&��Hu.��ؘC�$j9
�2U\)�*95}���&��o$��{+Y�W�9�,�%2�`r�L㚛 $U�
p�"R>}��Q�(�ߋ&�k�����Æ�C�K������>�D��*dX�Z��s�O�q�����;���rJ��m�p]{�$���΃"a�*�z�cg��D��!��:H���t�P��M5%�D ��L
^�#\e��ѽ�R3x.LGGA���U�p�Y�[+����K����!�Ά
	H�qc58@H�sLk�h�w�,t7㾟T-k��w������%$�ZwA�/ӗNK�{�i��щÌ��$i��>���)��w�:��=oSs{,�£_)�/���Γ��*��k! �E�T� 6�����T�&r�`I���˛�# ��ըI�"�~Qw�,|���t�C
@_C��:��|(��V�`�8�f�`O��`�?�G@/�0ƥآ�X}�|F?vj=����^�t�����~xv��j��1P1"�ӱs(�C[��W��m�_�QNH>w!Gp5ӵ$D�/bB��?�!�|n�T��RF�d�+��7(v�w�6YX����{>0����7:����c=hTP8�^����F��N�m�H$�D4���܇�2���66�߯�+o�����͋�')�Je"@v�L4��p>�����:T�6s��.]=HV;ޕ��*	6��I�c'�e�$�8N&~�A'�=��u3b,D��pb�dY��O(�J��"'¥б��wv�����/��!�1!����K���`�*������BC�;;;��8�02���L��B���1Q��@.'��MMVL�i�*eHs�;e�z�oX(���w�-)V��`�oÝSq�S�^��:�p�X��Ռ��-'�e�溛��l�r�x|��=��p���G��{ͭ��I��|lCCG�0 h%�>8�K��e�]\�͏���ү([�*������7�e�w�Ĥ�öJO���%���d�*2H�Ȃ  5�Q��Фu�5��2)��c��К����Wf�1*����nA�YapJ��ئ���ɽ����&j�ͽ&dЩ��p��I;��I\VU�3r�a��J�&�3�I������w����Ӟ��Ƀ�4�E��yap�L9�m�;��A[���$�8V��˛�*��5�!,�)�X��&�VP�g��>�ӗhܛI{��;a�rP��� ���2�2�EnK��O
����/���x�d	�#P�S~ą���k�D���?���do*�|Sƛ��'�	���
iw�u&I��
�ѧ��*5��M�����a�ȷWVvkSa�"�O������2J�gk����B����˯�.�oe�h��[}��٧�.��<������ kD~)��
�����g�`�5	Xtrg��7��������?�*���6�����ԍ���>�VUA��"���K�R��r�Ip�ߛ���mѶ
�8��bqt��D3� 	���4Ữ�-�
�z�Y�%^#�v�9�sj�f���%km�P1Sˢ2K

�N�0�"�9씷.Gc�P\�-Ѹ�d��"��i͞=�i�d`~Ӂ!���e!�٤{��aw�2��� ��N��=�O
A�1h;��#LS�����\p������(ԝ���g�M�v��z���N%	�뢤 ��~"���:\�&��ը�5I�1DX��q/��%�����K0��|/hmb�~6W͹{��{���p�,�H���q�ٕR�w�K�OA�xB%g����R�>M��(pȃ�R�B�K)�g�����{���'M�ei�M�A/B�f<J�<J��m�]>b#pZ�!#����ܷ�%��"���@�4����U9����0���P^		��s|��^\���������ߥn��F���b,���� ����d+�{o��"Xl�BoQ���h@ZP����� �pff|���=�ع��5k�S�3��3�'4m�If߹�}<@"�~>ww�00�1�rO���S��>=^��9���D ������
d����Ԫ�C���3w~����|e�*r�1���9``x��mFg�\�iA�n��)��&�\�ڟ}�-���v�M�N���b�Ц�{��-Ӡ���-I]�(���y�o�1Cܵ�qy:uǤS9Jr�!��C*ŧ��.dȚ�����a_3����2�� ]��*�����h3�lS�`�`�Q��sNLB��$��z#�~�s6q�a+Z����� $ei����*3hGV	B9RNHJ�Cw8���^Ȝ�� �w�u@��j��&M��ѳ���pG"�����ϥ͚�Y4:��p�o�J�E:�rY�4<�$��ݹy?� 2�*2i�[�e�$q��J�$w��[�\dͅ2��f|%�)���H|�,��추��}�9��ս�NJy	�=��:V�9@�&chϕ�EL-Rb ��Ms$B�˙?��P&}��P|-�j� @v� �H��M��7�d!
x�Y�S&L2)�I�r���hpb���{a�I��|��Y�k�^��
��ۻ�%\��j�<�!x�ߩ��'�[P�?ޢ���9����Ѱԁ�{�4jPٿH�.�S��I�%��]t�"`�i��;�6�>��g �[���ʢ|G�fAp��ئ�u�tA�2I�:�PJ���3�,��͆��1���#0f���~��*�X��G �v��c�z(<�C9�&O`	�?ׂ��=d�ٺ����F����r(h{[��Hԃ �zx;\��)ʺ��o��n�M�k:?@�!�c%dո�
&��M��6Gʹ^�Ƕ�c�m�?�i݄&<�N��'R�_k�_�@�:~�����QA��{BeF�t�e|��̤}.m���5����ʡ���c�n��T��^�?��ѐ3���"6��7i���̃��5�?U�C3h�-5ݗs;����̆D-�r��ѭ�S�_$�aTpD�c�63��N	���WZb�zG�!�r�#����.�#�{+'�&���Ğ��A���׼9��G���'ό���T�Hh�Y�U���n����Bv�ԔJ�r�����Ԍ;g�>��3���?��jI����Aj�b�T)���,{�fr�?U�Q�0�*_i���9}?S�[��n�3�evU5�29�� {M�qH�l��F�ѩ��pn���n�=pJ�#��2���/{�ހ�ɟ�-��&�X�@�(;�C��D�&�Ѻ�nkT|����Gݧ���ly ���՛��U�
ۇ�l=
S�S�,lqm���wA�Tp��i����j���'��rP4� 9s��M�� �k|�U#J���]BB:��$��,Z�?�]r�E�JI���Ͳ1���&��>�����B�D�Af�G$ M@"ܴ��&l�b����=h3:����p�w�B����x�x��92@��� ��9~�i ��T�\E�l©��[��kιr�T����V������ߎ�;mm�eY �z����`�_��N��9,<��lتt��1�zjzň�|(��\���.;�(�*���4�d)��g��z����o�f��u8�J@(V��������{`XA��"�gz��B�&p��:�F���V�[߉e�:=�����%OO���3�>�at�ڳ���>��]Pꘈ���,E�1}�P~��5��SK
�}�p�8���v�n-􀱻�7!=V��ͶJ���VZs�6�F�kF��'J��)�@7�� ����ݦsy��ׂ3}{����n�9�������U�vg7�k�< �j���Í-�`\RӀ��;��a�u^')��NB$"�K���*]B� g��4Gd(��d�������M�4��[m�e����+4�7�-��L5)�:-O웂����p�''Ѐ�C$�M�����p'�0����r�?޷�����Z�AR�� �
H$��!���̜n�_uғ
�|�S�zO���1����n���ڂhԡF�^t���Ϧ����Up�t��g&X�� K(��zE)� ��alV�I����d�\��j��$��V� Z؎󎎏�?�x�05���fWj�#����O�_Mڋ�� Q��R��~3y[)���ځ�յ��@���ho����_<r����Dp�MS�oɝ51��xÖ�:�J�Ts�����`/���t�Ml����p������
��{��2e��R� 
�~E8�ƅ��i�v2��kh�Y�`�'��#�z]"`��$�N�n��u�M0���5J>$���� 9���0.��P%����K��Y��T5�g� x����"V��)������6m��n�X�z�\�@
%dWzŗK�m���L�k�T<�@����5U�z��:�*��+��c�Sf���k�������PdM����(�cǇ:Du�x�_ �_<"�<A��^���m��"7D�t�.��9ǭ� ��e�fQ[�^]Ȼ߫*r>U��%�d�iԣ�?P]y�Al�5����(����-#����}&t1 `/U<�1���C�|�qK�b��VX%�U��5��ѕ6ˢh3Rf�
��2��z)�zD˄�����P�<x��E2D��f��7FZ�c�Љ�#T�J��vi��f���������	���y�=��Qv�@r #�qFqS4����͜�4��$w ׸|��N��h75H���:�GI�8[Tv��p�g
�_�Ƹ�Tp x	�c��h�y�dǥ�*��L7��µ��=Оg�C[2[�~�����7`) ��Wp3�c=ɕ)��%��z�+ '�x�����8���D�.5܀�W�y�6��W����֔��O���S����R_�Kؙn�ưJ��%Ĝ�20�d���H�b8}�%gu��5b�"PD��'���O桡������w�*�qʶ?ÚV�RX��H�E��kof'�SR���<ԥ�<�[ y��&�W̝��>ʥ9]6�~�Nٞ�r?��WJ����aZcO�ng.M�F��֤�J2�RM�����qCV��F���c?��WOq�c�Z�e��<��s��]�3��ܮ�:�+Uc��1EӀ::�?&z����b!M�Y�C�$z{����̨wΙ�WZ��qu(�������l�5�]���3�c<<{��Hcy2�����sg8�~&AKъC��C?��E���ࡖ���ZL �D�R�F����C.wzY\T=雵�O�l�!u�
��e�~��伳�� {Ƿ@�O�G&ږ�V1:qfʵ�D�Oq����g��^�h�̭��f����+[�f��X�� �C��n*��ѝ�-�6�U�%��!E$g[ߧ��p�`�SC-�~�-���ț_X/_�tx��D�x��b���z�´_���3�I";q�q����R�_�tpeggP@;H����g�֫ �N�4�������(�t�D��X=����zH-��Ъ�&��~Ѓ�����2����s������1H^05rͻ��0�^
}��.�~ƌ�%v�V���EhsK߳��s�xӕ!K�I�Piϱ���E?E�AGX�#W�Ҳ������!Ẹyv��UX��'�#I�qe�ރ ��J#�$˽;�4n=B�M�f�W�xޱ��S���.���� IM󰤣Ϋޕ�wLf��+����� uȕ���r�d֭ȟ����^ P\�#���e)�mR�AySa�7t�H�A�L�-�Xي��bE��x�  �	e��=f�z R���	ߋ}��#�$�[ ݴ}�b��1�|t'$�m�W}c�uXl���>������i��j�[?�Z�X���X�������&Lac�g��Ķ��u�a���|<5m[㍼x���E�afoȱYw٠V;a� �?�]�^�8J!I�pTpa <o�+� m��do��:�P���Rt� v�E<E;q���Qх~& ��e��1�DH�y���X�!#�{+izA�u{��mk�c��#T��R&���$Y'���P�J4�k�rU����E�Z� �x+�=��5%AW!�_�q�4t�r=$�Y���t��5�(�y(n}	꭭�SfZ��6�ʚNhH��`�V^��}����`@��	<����> W?�:����J��{Yotjs����b68:��p�R��+鼖���FD�z�:�?�J�>�q`P��m�0��-ߋ�~�X��w�$^�L������$wk���$�T��y�7n�ܠ��g�Fj��s�T��`�� (U���_��4;����#3�,���Q�u	���q��3��sO~'�u؟���)�'�i-�N��a�� '�ޅAW��@ilb�>��8ٵ�T˱��t.��<����]�m�0��>�I�M|��W�5�S@t F�R�)
���Vg��y1�:enq��Q.[��Y�P0ǟ�AY�6U�i�@�J����9�
� @<�ޥm)����A$��^��5�G�K犯w�f��ʐ�@�&�H`�-�{R��ޞt�,0Y�� W �Lo�C�?�Am�i������l��+�y���JP��nj,4xZ���q\G�^j4!���H� �73�6P�UO�����
U�>@!ͱWa �JL@���q+�_6d|�x�g`!���c,#b��0F���^�d5�p��l`��̓�0��\W`1aWQi�\-E�Xc�ҟ�KΦ6��E��
��H�#nNR6	`���#4o�}�(�N��|'��ٶ�d-:B}54~\�Pn�g�V��\-	?u��˭���J��=�-������f��U�-:4�lx)$WN�&�����Rƴ^d�6�6h1�/0�p�#�r@ImB�-ԩlmD�lI�����N�����۴���`ľ�F�bW (GC�B+y&"r�����-hN�=�� ����/�u�5�2{�3n>�r��rQf�W��&���
.4Y5n/��_|��&�^�
�N�K`�ȱ��_�]�N��?�
B��s��=ɭV���� ��(�f^p2���}ǍS�
��T��ؔ�<�kX�5�;L����I�_^�.���y�ܑd~�Pc��y�11k7��7�:R��A�B�ˮ O�ݙ41���#��p.m3Y�P�R:W�[&S�>>�jS0 ��h�}�݁{~/k�%�h@�S��r�B,)�;j�ښH�� �_�N{�4�S#�R!��F�}��d�P�������vД��2�Ew滲-��.l��9���9p
jЂw>�8�E[��r�5�K��Vg�vOy�v6�J�,���X�+��:�V�����ͧB�(�A=�ߊ<�V�h{}�J�����zw&�Ԩ�-R��IS��Ky#��@m���M����C.�מ8���b8�V%� .0��]�%*4ot�K��N���p��Y�E��z��EL��yG'�ۣs����J	�͖��K�͚	�9�()����f���
����7�����潣n*�sx^�D����S�q�_���|p����������C���b�c����Zh����kZ�/������;j`�5�Τ���/́�:'���\�T�naCݨ������]���݀��Ш� ��4m!��)��J�?�q��1Xt���۝�7|�R)+N��|��.k��w���uahk}�8 ��o��H�5u  �s%���d�n��3��qe`��s�;����	g��{�'��!p��f�|2���,�F�}��ӄ"?�b/��9��u�?��xF�x|�۩�\����k]Ŕ��#�'/.tJ9���o�w�m_��:+*�Z�ڨj��w3nJ�
�����ް��>s�ӹi�Qs]#t>�֡h�V~V�Ύ����J�C3���,�P�5Vc��ۻ�B�+;�K�nwh�Z MK�+a9�ղ�Tܘ��{�~�����ߧ�T�;���-�m���&1R 1�Еo*4^�¼;!���x���-�>[K�B�#���L֢���[uO�3�?��~O+�\R��,&4�� ��ky���t�=��h}��}晊�ɞ�R�*��RE]�2�:�x���4�
ͭ�k�x����v3\����U�+�GTH��_VO%�~�-
ֱL/^^1{�d^���T%�˥�|��
�ZYh�\�<?�1^��c�E�D�C�Y�P�5��/Ȱ��(�}��TSJ�%P�=s�Ȭ�>C?���_(9D��>ܩ��#��a�Xލ-#��:��d���F���E�M�(.UѺ2�#�`�R{�t���u%����j�]	LS�B]z���-�Mp���~����k i�'�(�>�ixW��%�y߸Ew��;��X�߫������3��"a_����d �r��!��?i"�r���PA˭�$�X��4Q/4|a�n>�p�O��z( f|M	��#+z������X���z� �u��8`�!z��|ʞ:6��K��l^X���Xh�n�gi�_��I�GR�0��{u�!uCϱN���tV	Z/��-��.�o`�B�E����U���ec1r�ҞW�?_E�>7��� ��F�l�vF�=Վ�F���9�B�����	6���}fĞ�%L�򴒆�jϑP�ę���ޏ����� ����Xd�rV�404t)O��dӜ�è{��%�ʍ'_X���t����؉2[v7�o�U�F�aX/>��:n��:�2�y�9�.���5�;�<5o*�ӕ"��S�)��Дq͙D�tw��R(GS�����$��8%*�!����^G�ɾ�
��6����9�6��{�5��`��w��T�4$Ò�9��_$\�i63+�V���A�v�-K�>o�������T�\ڻI�@o��&�B�gW��V���+3�a�W�l�WQ�/�.�ڦj��X�)�%��6�����ܖ�ә�m+ʾ����xXQʣh,掊_`�KI�c��̱�Z3�~v}ʴ��O�����=�Ŭ�[ؑ���譄֌���^���SZ�������<+���	����og�����1����Jy/�^6�R�o�j���`��n�s;���{z[(ә,wzZ,G�c�(�=�YJ
�k��zph���T������N�ZD�m�\�ӱ`u�b',�����K��%�$�,F�w/𸴵�-�f>���WS��>6`+Z#\3����J��I����am7��K⼣��^�k)�pF���G��`t%���d*z՗W�!(�,��N-g�+��e�L�ٜB��9ᛸL�Vie��-�&z�����f��ѓ ��LU�N��bh�T�Y�k핲���+C�U��0?�'�!r<pW�c"P
-��Ni��Ḝ�����%`ŝzt%���H��2nhz���d��Ħ��QИbpSG����3�q��v՞�����\��.�T0+GKcb&��pw�S�N:U6���x��2V�0�^�A��h�Y(	|G�$& ��5�`ҦSH�	�#�	1��E�)�L ���X�E�������>s%��h�<,�Q�������V�>*�y[�ל��&��~4�ՠ����g�q���ϕ(o5$�Rb`�׃XЖ�4<�0�ٰ���4��@�T�I��Ř�eq�>g͝_�:?��k�9|�.-m�9����.�1�R��í\ѽD��z�L0G2z[шo1}IA�����,O�T �*�}RñFQ�M�������F�Wriʩ��ǝ��݈�P��̝�LA@k�SE��i�G{�aakj<�ê�h���S���`���)VS3}�R󰾺�1^���� '��j��7�bMx$
���c����oڰ�B[�U��Y�~�$TO���:
=��Ҝb�'�oT9g�g�Z��GD�q�7"�I%�Y���l9H$���+�]+B鲥�gjx���6ԙ�*�.����|r>�(�V'f��T��R�ĺi-d�,p��feP�wI��l�"��@��yV�m�yS�Ȱ�s?PRHܛ��kg]o� VIe�jl�)1�J]6}V|)��,<DŃ�&�h4�C�:�h
GK �:@g	<Iў���F��xj<�3���K#�7)Ӵ�	Y��O/<"�x�am�v��e��Q,�Xp���S�.�9�������%Z�Q��"B�r��sx���*�t�!�:%�)Psgx��A_�����^n������J0����7�W̣,B�W����̝[�/���/P<�+�	H��������u^�y��Jg�Ȋ�;}q%߫D�܁V(�TN$��z�\�{Lx.98���]�=|����C���2"��$�"TiI��Gj3]R����H��:)����%O���u����ѝ)�f���#Ո���\�p6r�2<!
i�d�������i�@z!����bzw��y���X�oXt�lCE�.C�Ԙ�Ĵ�t�e�w��ѝ����PTL�I�[Q��ьt 1�g�yF���ˉ�h��>/�N�2�*k��C*��Z+���C�OOȫP_m�?��B�rW�(Ժ^ײz���F�����r:�*��]��ϩ�	�'`�_������[]f�E��w��vv�U�R#ǻ,kiǰuM�
�an�D�+F�S��<)�]6�����#e{-D!5�i��Z�E���b(ӽN�����.�_�\�,w��Vr�o�� Żb�[��3m��H���`��Z������u:1?-���%�������qF;�nM��yg��2�c܁��m:	�d��__�P�^m2��4�L�2����x�]�^���+�v��^�� �@$�k��2��@U$o`��˘�	K��O�֐�s�Q�W�Va�.x��<}^6���@jG�x�N��x����A'��KM��"�VF!�e��|���f\u��.��(�K^6.��c��x�J=).6�1
�x�z��,p>�<m4�dt��9��a�&"�n�od`99*�o�ݏ�Y��[<xhN�������9<6m���)�my�NH� )���c�y���Tnus��J$r��B��3��~T����I,0M
6pwM�`�˞AM��欥��N��^�s!�)��C��pZ!ڕ��1	�M�7@9�3��k�M�Ba�+e��i��9�-&���"(�=��˨6�N�lMQT�cs���#�iXk��QQ�8I_��d9w�80��?������Y˧�3�>�3,��4^Ԡ'r��Z�WFzr��|���q�F�O��Ou��n��1Za��N����\����cf���y�;|��d����v"B�~��ؘ�>�<Hg5��ի 5x���1:.�x�S�����l�a[��|S��/��[��hH�!X�
 7����A��Ӹ�.9>i�],ם�?m:�56�V�jaA�<��n#��S&(aS����}2$����Gw�1�{��^"�Vi�!�%��������H�A�Q6(u5��>���9B�}���:��l��̼�fyrD+}�ۑ���)ݚ_Y(-R��i^��ǹJ7��h���%�H�L�?��,=��|�.��ȱ�ez�$û�T�B0M�g�V}Vh%� !��qf��%jwǥ�r�[9���
��L*�Ŵ��������]K+l4/�D��_���dN��=��Rc�\����xV��Z�Ra��ߜ�.b�+��t�����[ݚ�^"�Q�Bކ���g�e�>��[��d4]Dk�)����X8��xv��o}`��^pϹgt��G�e�!ә��NgG؊��eI�ʝ$Z�qZ���k�7$kh;��(��m`	��\���8��H7��6d��	���rw�\���/��~�����6��>��9s���1pB��j�r3BW�;�bò���^���5��9�.�3U��!�����x�|���^���?�j�4*�I�8>�k��摚F֭c�����F���-*;�����j�s����7N�	�	�@,�M��Ŝ'C��η-F {|��иEk�I��Y\~Br�l,@~e?u�]�V��ٝ��3߹���Ic�kF�FD�z×�|���O[K��Q�X���t��s���[���1տ]�N�ki(�n�ւ��o����
��Ϝb�E)Ե�i&8�|�����}יͯ�����~4W���q�eow�憌z�ޢK�3_��񧨭R��<��l��V�!#���Q���R�U_�D�����5�0&;��=�<kG������l�e���p��΁F���<E�;~�SE�i���S�z�=�f����4?H(\���\�_�o����*��좬xڞJ��������{OH���Ɉ��	�e��|��	�͜5yZ��7m�?����'�E;��d�>AR�T�uqZ%-o�����M��/>qOa��%���V��W^�ҍx�k�(J��y�qˌ$#��k��R�L1���&���,�e�ٯG��T�4^}A�f:2��
h۪0��]3��m�c�����[���a��dT�Z��y�������^5�EUfr����'�J>���	�T�ڞ7F�ǆ#]ɲ;UB�F<����b����Z�nF�巐,����F|��?�����__��aҁ�R};Ƣn軆��t1��fDl*}����֟w���)Y�����{6:�;�Ȑ���w�1����c�z�?�_d9�d_�5�H���Ύ�N!������*M/d�LA�T��<JuxF�P�r�PQ��/'z��>�m.x��4���rՁ����[�eR6w��ʛMډ��;���w�7<��S�<�\\zJ�&{ǡO�������/�z} I����}��C�zшL��5+���}�<�F��m���P,l[�{헑�O�0���.�9�$�Sp��=�k?��Yoŝ �� EÅ��S��X�̀���͆'�6���ƌ�]�������Z7�����Y��ܦq��_�}�j�s��7��3����8�>���~�h��	=�,�CcU�}�O���+#Vp��8ա�MN�AW��k`׸��{*vXؠ�Zpv*Oi�߉�O)݈����@};'-z6<d�ڴ���
�o���r���ڭn������i�j��\�/���=׌�W[.A�d^(�E������[����ڣT���~�y���T0�O gI�h��-�KN?a�	�|A�Ghwk��M���N�7���l�P?P_�����#z�\?�Zf�NR�3���{����;hh�!�3����� {�Ks4��[X;������V����<y�$�w=u:L���̇�������A����~J�ޙ��糎�c_�,wj-+ls�c�=`��L�oKsi��"�x�ݻ�v�@d���F�3sv�B���S9J|Ď�E�5���,<!pE�\H�U1̥=����2��1��ma��Z����~¥!*�Jb�2�:�e����4�����a'�N��8et�K��K�p4�c�@Z�l�����~�*����3�tF:����"Q�_����}'�������~:9�P�=��D����d�O�M��C֥�vZ,�\���|r��Mn�ڙ�!	�z��󒇁r92Ux�1n�m�8_t������ʹ�@	��d�'�;P���2/r
�/�EE��~X�Y���m�8�g�`X7�c|���_ڤ֩���$�H�aа{j�����F�4_�NG
���]g��e�wq��8^�C�]���4��i:T05)U��U��O��=��H%4��t�!����S�Cή�sU_�܈� �a�w�kc5OE�ʹ�<�%���
�����}�z���z/(u�Q�گ��^�חp�ԏ-M�p~������J���x�����]��w�'+%�U�0�?�jU3s���CQ�h�g�&��̎L�J�bS����@Ce����Ye�E��F��G��U����1L�Ѷi@�^��p��������o��3�h 8�zȓ��oވgtT+#���v��@����+��A��i��3_�@�Q(�v����Ѫ1�����W\:��Q�Uo�9��v�W�U����K��rVł���t�tW;�՞�ʝD4ML�A9��J��s)��%w�Â~p�̝�3}Y��ހ�EY����wG��~���,���3��	��v��i�D��GN��B��!��U>��od��[���	�����m���6��~����h����Te5.j�9��XP���G��U���Р.�6����5p">�� a|��-F�1���s*Ӡ�YA��АW{U(��|i���'����?�'u*�
boaI������?�/A���{q�Q� 6��*uҿ���J0���4�2�riSşm�Mʾ�?tNuL��E1x>y�/��X�3�P�|>��?��K<̸>�m�r��a�<O?���$��M�D���l%���#�[F�)k�2g&���<�7:�p��u�Va<��� �	����&�tb��m
���m6���Óuv��Jq��� ��y��c
������!B��>@��I�H�ܖ��b<EmG]�i���^`�#��Ǐ���|3�DU�G�Te��s{�g������q�O�D�����]rmr��Hㆿ[T�ȁW�cQx4�;<����&�Ᲊ�!.��O{�\����ʸ�o}R��B������g0�;?�pR��K���aD����	*ǣF�l�E�e�������#�Ӫr���dP��e���ϱ�@��z��z�K����W2u�}`{�F£�6T�ڈ�ZU��GlR���̊�0���y��XH?��m*|��x�^�7�D�_�#�/���Ar��A�_���I�k�W����S��N	�[on�����?�ϒ�c��n(U_3�3r��M��̽�S�{jw��Q,�<9K3�M��ڞ�]����F�m�ork�x����{ӔX8	Eڤ��D�����z��0MJ�~����}���̽�U拆����S���N���V����{�,�%��{��G��'����Ny3$����R?��������a����X~GP��;R��s���J���!��kg�&5ǡw�<�`���o�v�'s���5���k�P�~� �;םS�>�0\�����DL��Up�/��Q��=����%���D����������˚���}.;��w�\�	ioЭ:��v�+�"1��`�\+;��|��m�D�f�gѷ'	ܢ���Z/�[ c�"t��c.��;���S�k��4<t�$y�1>G�%���Qr�{ȢylIz�-E�?G	���k���(g���Eh�TC��/GP�l�3��P{9��9������>�e��ƿ�:�����'����O�$چs#�ی})�%���Lf�$>���03<�v��mK��>��>GU�(��Ak�ڧ��O��X8�D��!m�l���1z��:�H9�-L����0x�w�o�qG$�*:�Z_�x�7�K�J���t/\��B���wi�&]�$����pu�
���s	DHY���R��d$�[F�j˛�0�x�F<���7W$�ä|�X0�͂m�ˏ��qG̻���iE8}�����`����9o�q��3_�|(U�*�օ�(3�Mn���"��g�V�֤A�$�ݨn�v�穅�9�Z��g|ޜ�x��Vy����l�����ُ�d^�e��F�/8��J�n���l���'�0�3uv܂�Rm1eLW���>SQZO�4(9�;�ֿM���M����'�d򟐩��7��_'���+��.S����9�x�����sQ�.e橿���d�yJwI>�pXs��PC�aǫ���2����E+����$��J��㳫����Wv�Xt$ݡ������Z׮y��5<R�x�ɟC�WW�ܐ�Zƨ)İ�(k�k	Lu���Fi����p��d��ɠ������M(��]�#r�~SM��	L��E�y���
ZKi�A��9~z�}��;D! ɛ�{�����ޕ��.U�2�ԯ0ye����8\�,l^8[���1�{��"��J�/9��"��"�\'�m��&1L��9�<��
(G�q\��`E���s���P�:T�zx�W�+¬~{`6�A��4؟���qM.��5o@/E7١j-�T;[�&�q�-�Ak�͟�C����Ó91�`���c}�FP�Z�^m���4�v����d�iQI}�z���ÿ��C�!�y_��/�V]�/�=nJ�n���)=�؂�R�^��W�x�F9z��s�l?`�U_Ӡ�|��?�U:D� ��@��{����%g!<Q�A�����j2aT�!Zf̑��y1��6��25I��B|M��4Xfb��M�9�h{}J��t
}>���1X�	E�!��Ft"��Wx=����I;�U��jy�h�.�|�
���;k�;��5R׬�����.���v���������_�$�~�yf�J�^�S���5�W��Nf�S��/_/.+cNMM�4�h�����q��"�������e�k�[@��MS�Tn��I�*)*�|��,~r��+���_��si)x�Z[[+q@�U�E����wFc�C͉ol�T���ȅ/%�(r���87.))i���쌳h�o/������C�e�3K��щaFy@X�֪q;���џ�F���ˆ+Gw>�������fgei��q蠩l�pΔH&r�������B������A�v��I�A_��,&+#�aw�hq�t�y�=�9B�؂���������N��N(�{�ʘ������v���%�;���эV�u��q�<�m��4���2`;�f�x�䅠�)�[�Ȓ�J��KtOq�f�N��?:.��K�!��U?U`u��E�p�s5��Gˇ�.Ec��Ԥ�O����4��)W��(�+`Z�����i��V�U�C��vx@k��b�M#I�{L����!�A��h�l��:ʣC��5��[�=X�)&ٯ��A���1<v�����+x���Ge,w~ �F��Sf>����"�o[���jB�z�|V�|�����wHC�?�-�	.���+�����e�HђKz��?����w��d�R��zG �#mk"�v��'͛�.\GPA���#�?��v���sL���� u��թc�@//�w�!�b�n�#S�����u*��'�|�X5��+Z��;�^-�h1S��%��B`�.B�!�{�Fd7l��=�S"!. 0�1��/	�0��&ɑ�䬓+�WN���'p��|-6�+mT��WA��[����و�Έ���q�O%)�$�ڑ*&0�/�F ��h� �rLN\���U1~;b�y+M���wD�T���i��y����u��WP |���� �R�I�Nj1"��ыk���X�:SGt��{a0ó������OLZ,�iz��D_�O��'52�l���td"
x���������~����)��@���(:��#�D���B�����3�t( fF' !"핂Ҫ스Up��:5( �� ���q�v�oc�Q7'q8�T]r��	/p,q�!9J��hը����3F�w iP���D2��F��x�<D�),i�,�����՚�͎Et�M�԰0.>t�`�u��O����0�����/tP�6�o����ԩT�N�����-�.��hB��kt�вګp�7FI��ź� �����~��u�h�<�34T�B�������:�>׼���UG'�3�- �Y�F�����?N?y�D�����b�j`�V[5梌��A�K����ccJN�O�݊��mO?k��Zs�i�g�M~��v�G���DA��(T!�N�#:K>��8(�鮁�lk6{r4���#�4�J�|�=?�Z%߾]�-cZĠ	hߑLEZ�h[�AI��T��0�Ù���NM8�N&��nу�O��2Euy����uT�J�i�Sj٠�s� ��J�㥞��	�Ng�/�}K�n��)�99�W{⟓�M��ݯDl� U{��&~���Z� ��(���ǜK��?���o�e3�=1�<&r��jaKgEÜ�.�a�o����Pz�|h4r꧀���0go*ʺl'�F �ڋ8"x���k�o��*���z��� �p�9]V�f.1Ul�Q���^X�h������U�2����
vS?��U��5Y��eu(=&�o��g����TGB�T��6�_�)*!��
� �sٔ���������'y*G��Y�A���P"�@,��/�yD����J����q�$��+c�+%E�ȱ�hgr�4$R~�KS�����*��� ���Eʕ>��H�Ne�f�g}����r�ؘ��ġ�{�b���a.�վbXH^ X��)�#.�kXnL��e)@�.Fr�,��+�JɎ퓉�eA TوJ���d��	]2.����(��c>� ��1�܄�7P /xY�IT�U��=O��L�\���}���O諾�XYpUޔ��j���W��w����.B 8gg�N?9V���G�1�W7�~đ�s��	�%���b�~���OG=����V���+�h���9�<�^l�V^��1Έ0UL�x���5f��������O����5������χy�HH���7�b�X5N��<�:�YYu��i�������Y��jsǓ���}�!Y�3�.l�@xSP�?���g����9�ޕpw �,�(�Tj�V�+DSk,-@��х����D�<ԕ�lI_�$���dBJ`+��a|T�v_���t	T�_�n9OQ�5��=t�<�,x\j}
i��\����4��F`Z�Ӛ��â����x��sT�p�*��	Siv���$�]�v�G����X�Gp��^�w� e�9��q����w���Gv�ǟ���qM��|P��RR4��pJ��	y4"��s�(�2���1��	�Ikh�(�A��s���>��FH�_�g��������ѷ_42I�Dw�H��x0m�9�kK_��4�\���!���Sx�s�]\�}@�4��7W������6�����D`1|�����Q8�%�>8F�)wcr�hk����:n��M�tI�	3M�3�t{')�t�z��V�	3�[VM��̴y���)8���#a�G�i�6r'�}1Z-YhIv�4�}��a������'ێ��O�<�G�f�b�c�
�K����k��<8�����~E�����'��Ø!'/�w�4kq�Q\K{�ر�W��i��/��(=$̍W�Y��נ���1�$���?�!`޽av��w_܉�զhF�1b���O)�E�P��<^�(��͎���*�x����7C!u�c�ku}�$��_�r����
�Q�-��������2�#fk~���z��g{����^�0[}<�� �_zu��n��9&�Y�q엤�#�/l�}�4��/�G&^ׁ�4���}��vb�z�X�߿�\�l�2]I�T$��C�O�O(�����-��ᖍ�����A�-���m��=�ֽ��E��!A�W{׏G�v���)�O�����~��l�u�_<'��8�յ(5i�ْ��^��.R�Get��^;a!��p/BBs�;�9���'�>ۃ�m@�i)NDY�QwEb]^�W}�ŝ���-L�G5a�[��gy�����}Gb5����'1�x!���C�$���c�4���M.(����u��#ǗIᴮ�k�����	ۣ��C=��'�T+$@�h��l�?���DS���G�`����_�,"_�$�jձ��8&��q�%�Q��Ɲ@�H٤����ax�ջἂA��Y\�$ZL&��)����` ��Y�ɍ�V��>���^��Ͼ�>(�4���3,�
7�<vp��0v�yp��(E#��]�lBu����3�h�#	'�r��m|�}LԹ��P�ҫ����u	������+3όc�{P�� �������/�Q�$U¥�/2���|nd{'��ـ��BM��`��oI/5���^��֓6�$T
�=�r@t�Zh��tM)K�{��]�*wo�#+�@/&��I�нNu�?"dw�UP-Xhf�������;X����Ŭ3�B���q`���	��)f[���҄R-�����2D�U�-y�7�z��<����IQ-�u�rY�������|M�E���A�D�0�&Н����p!2�M�W�2��km��Z ;XK����"HC���|�n��ˤ^n��Y�n��I�jڥ�au����I�&����B`����N2�vZ�����������(��L�J���Ȭ�Z�T��{��=��G�ӄ�Õ�~��e��[@�K�0-6AU�l8s�쑪�'���:������j֎{�Bڰu%�����"�w �P�[ʅ̨�`!b����ӿ�r<�G|�;>��z��'��$��ًT�#jT�·��S�1[��k���Lf�O���\m��ғ�;��|&��5�^���l?��mA��wd�V�"�K�"���'����BY�HF#���]QW��h��z�s�bq"�Gt��h��R��z��V��IoQ�!6����Z"��|�=��Bt�y���ҁ0���������#�/��R�(���7�/{��hn�+�
�k�zB0�Bh�;�=�\<� �Y�/����Z��LJ�ƨ:%~xv[힨��]���«��8x#l?��gߘ�0N�KMr���u��_������ZԴ}-���N40R�_�`��o"�� �Z��3B��Oj��M��:�.��(:�E��]���2�>,�^�ޏ��T ��ċ?��!��Ȏk��Bc�ф./�J���r;�Q����|Gd�)���)�-l��4��xf{�)G��;H�@�9�BS��QL��� _)�?�����t�i�e��q�4<Q�Hy����?`�<<��gUP(<�NY��F�_B����|�y�J-y3�q�W�"�O2Ǔe��z
wn�B�Tgc�e�q*���u&���7��!x��'"�c?�e����ۈ9܂-����6��u�^Q:�q]cl��+�B�.�f( �hW���_��ی���O��9Pe�[)���c
�}[/�Z��ӟD�B�p-�M}﬎@>�u��3��a�&�蝔�S��mxgn�y�m�%dE�7����-�ޯF����8�s��׏��o�K�V� gs�-w�p�'C�8?}�<��o��_ș���D<rI���o~㵎��h� n�z��-w7sӨ^�{yb��9��}��$�˘O^���F�J�#�ɂ�E�4��n�6�~�_ ���5ۿՀ:��(�,�C�M��c<>���]�
"!� ��4�½"1��C�9��-��{��+��Mn��˝�}�c�ps�L�U E�h!%ቚ��qɣ]���X�+BQ_)�C�����[�`��:00N{"�O^�dB;Wq�\���q<��Ë\�EZ���w���Wi� "�0N�R�0�&��wq!���2��� '�7঑��?k<��؄��9l#�e��a$,`�A��9���PZ]9;������ �O�R�<���,h=>{ ,<7x�  ���g��A��2y��m�T�w3~�0x9�0��l����ʸ�8��ݖ~���AO���\_]ഘ>�7���I�����P�o���!���di�ʮd�ZRI�ʖ}ɾ˾���P�.���}�$E�}b0��`��`��9��<�������+Μs��}]������>G$��v�n�,>V������Vx��'�������
��~҆��)h1�'�d�w�1�Uq?
���\Q�n&�<''���2D���=K^R�<��Ot�޿�!+���k��o)����4lF9����b��@�i��H�r��T�?���\�騊�e�8NN�TI��E���������Q�x���S�~�j̑Qg�!��k�~�u�^��~��\ �;�5t)����*u��=�%�5�?!�|��z���q���dvQ�[5�撶�Q�K�E��s%S��j��dV������]�3�߱ݳ0����u+H���-I�.��h�V�"۝��&NP����DW�'���O�D���/`)����Ǡ��n'}���<�M�<8��	����?�8J��n����vD�!��� �@jlF��F�T-^-��a�T�bF0�5��x��ӿ*��~\�o��M}��|��L$6K������;��	�e�g����w��K(9Q�z� =�E��y ��`;�����a:r���&T���En���^�����)�k�P��%�
v-(}B�'F}�G~ȟ<& �j�_j��&.�R�M�2d*G�����Ɛ�6��?}��;���>�b�_ �(3�h��^�S�8�S?>���&_���/5�W�
}�sZ�8�9��/��s)��_��_���#h�HN6�PȔ��|n2P�q���&T��`��s���NOM�U��q��٫��e�.���>X��X%�&"�^�MB�� �{6��L���%�f�\���c�ŵNOB���^B�	�����{iQ����<�l��P��_�0��T���g8�O>��T3�R��a)��}�K#�m����+��#z�����4'3	�]�-��_�t-�{����M�E,��+��e`w��un������PI��������Y��u��?�n7�U��Km����?���~�-B����<���;�~�~����R�d��q��矣R��D>�$��ŐI��FȄ�I���p��}���~y�R�tt:�t�߄5������`�	ȟ訁2�wc��+�u���$�����I����������\����c;��\ur�mi����K�+����o7�w���,���c����0��^I!��n�M�����X�O8����	~�ء��.��PH��G� _���).-qLى�5ùLo�+��Q�%c#'�#ΰ��U7�Lw��s�I�L�Lղ�����7��aǯ~��r?Q�gS�5i|?�� �}y���z_��^=��F�p�)T�6��}tz+�K�)��g/@p��i�qB���8>��	P��:���	O.��ZT����2r�5���|����+�|��_��n��4h[�u�X�ϳ�n�폙�K��t�ݒ1�꾹�[2�tM��F�� $�)�jܯI�kR��Eg|Z��B#�3�o��7q#~z�}x�w.�9�ib����>�9��I��.�b����ۖ�Kx�O�RS]��Ķ}�`d�~��yV$��IP9�r��E�{/c��p��B	��Fdo% É���P�͇��y�bɄ�=2�`U*l��3���M&y��������j����NB�.g�f���ӛ٫ObH&%ނ������j�w��ÙͽD�>O^x� #Uև�5�d��V�71u��cK�����}�Xh��x���j��{�cp'u5��k��I1��ӛTG=��;�U�!��l�l���h�{s^P�L�Z��x�Ң~��I2�� �<�L��K�k�
��j�_"�!L�����-�D��	/��Ke�>gq
�l����!�l��#��g7�:�ҾT�zs�
c�u���Hmpa�4���d��o�yo���z�i���3x���?A@�x~9u�5�3�A�&�-�H'���v��8z���u�q��_e�?,c�>���R:+"���_&!��1+�bV�4�Ժl84>�l�x�~u���.+�/M����
�u�",�R��7���\���ׇk���oN�� o��p�ƠJ(M�䦠�_ek��]�bZ�#�j�Iˣ�̧���RG����q�4�7,T��ͭ-r�~\7`Pi��%8U���;�������P��Їn�#�r��<����؃kK���N����3�,�1cz�O�s^�y��4s�%[ՍKN̯�i�rHf�R��.�����jjj*�8����Y؏O���Q?�add�j������Z�U��B�~b);S�je��٘,-��Y�b����Ӯ�f-cۃ����đ������;�]�AUN��ܼ<k��b]A;��KnW��uE�n��O��o�����L=�%�94����uxտz,����O�X���c�$ hk�W}Z��[V���8�᳷���ݞˣl�o/~���_�o:s�1B��mD�Lƹ>�-����O"�Q貲��[�T����$�;����L�Y�E���l(�5pb���E�Q��@>u���-�Q�m_iAwz����̊t��Xc��	+��%�MF^��X��f���$�4�,� � ���(yR@e?/M�����c\�w?���ɢ333&�.\���.�n�@��8�([9�W�#��#�í+N��J/����'-��M�;����SC�4��a��N n./c�끦<���ۨV$��p�ȝ6���'�~��_>����{�p'��	�&C���5�������������	Q"T�0���궕�[%/�|Ge�N��P���k���t�����-���f��ne^�N{��8���r�T�T�z�h`p�zo�X�e[�͊!Fո���g��)�pR�sXC��R��SW�j�n��K������g���L���{n�6����}�qp��*E����/�El3��ҰgO�q�5��*�w��@Q6��wv��66-�����M���k� :�G��[_i*�P6�bx)y��<���\?˻���
��)	�`���j�d=Y����Ƣ�GtI�n�4�#ܝ7J%�jp��	a����w����g����:��XJ�T�ݜ!v{�B�q~<Fqo� :�+诋��9Τe^=����h ��^�'}y�%s�A�ӊ�l�����+������s������@<�b�K��L��Z�$����D�/=(F�{�e[d��PZ潅]2ɴ���477W޶|G "��݁\!8*)9���" �4�@`3�Ck�;����sK�<PDdޛ�ٛ��B�}"Yw��T�4Ҍ��3qI���d ڨxߦ���Y�#̀�xWPP�����&�_��y�Һ��A��#�x�SL��轝�Όr=�7�i��>��Oܙ�~��hi�q���DX���`�����C��·ӈ�zr�9�+�|�x6�4��]|ZN��A��5 #��/o�]��3D���_\�4`��9�G�8�h���厝c����l�!�?''%~��=4��6�n"�dм���r�-ߕ��)|-y��W�_!X5�� G���h�z/V�ge|b��;��GA�9��V�4���oye��W���c�X#�y-�tg�$v���i�ţ���o"/7��뺁�����L-�s��k�ѣr��Hn>U/p�C6xy3����mBh t�{�o)���Қ������]��5)�V(Z1���ty7�"E�fC���p33g2�O�0ۄH���8Z��B��/�(nX*zM�~Sj�۽��H�.je����oO:ל�_r0%���u,C�1u3{1\�⏌��h{����NН���L;�G�FV* wθ��I����$��;D�Us�^-�-����/�c�7'#EeX�8��:{��9�{HH�h��I�P�bS�+!!���@�x����}ܫ|SN���FA[Ӣ[!��!ؠ��� �7-�{k�X�y����� 	?a �r�"�:݇�}��K��T����RӗJ�c��H��}cz��k����}��M�b�x���E�j�3���Vf�c �|L����ݗn[K�*gW��Oȝ[#W����R|q�Rз���q+4��}�Ri���M�6ŽU�`X!���d��D+�mM'R򔁷&��	����5���o``�D����O��+����U��Upے$��h*�5�>���p"���Y�As�N�4,�n�'��;����:ޑ~$zj���kZ�1#7#K6kA��P~ Nܿ��W�UJ�"4,��Z_��꛱�_5l��7�nN}4����$��J��q@9q+�������͛d�?�Լ8�(��"��`��|����ؼ��a
e�2S�^̧�������$n���\�B���P��X�jӕ2>ՄP�uE�Υ�o��%S&z�D�qqj"[�����;�؝NӠ�HӝDI�B�h��*U��O����D�h���*���^�܀d�Vcގ:?kmU9M�a��Wy&�|���###��u�E�nI�X�4wvi��M	Zv(��,\R�`0�!Be4T���8�������lzF���%��e���s	�	Sp�%/L��-�`E�~FӾ<��� �����0c )ZH7��M�6<nɈ�rb(�id�Y�"r�/cOʷ���O*�8��醌ע~������ﱦoRR�w��c�z���B7�R8��1o�L� �w�;a��s�؇�Ur5���ߺEl%5��"����=b��V*`FJa�-sc�b-�&�����5����&>�x=_BW��C}�<���\��HB�Fp�_�D}�=I��/��Z~�:}'bё���|�wR]	�B��� ��mZ�,%�����a�Ґ'��D*�m���OE�V�'q˸���T����\�����&��QM�����кIic�rJ���M�yyn��*'�U�\_��X%�eߊi�}��m�?����[�t@8���~o3�@QG��h.��_6��7���oRӤh�����9��8Y�aո� _�A7�ͽ^1$��p<�O�W���ƌT�����څ��&͠�W�������mT7�Kn)2�4�l�ecOx�@  ��s�vm0�����I�Ҿk��o:H��5�����6��q�@�#ťi��4`Z��n����C�%EF������G�l�l']}��d���/�U}<�����cw��������U{\M�׿�~Y_�x2,�_𔋡�K񟝝VR��ԗ4m�{Ct�7 K#��uH�n�w�`4�l�]u��M�ai�޹:M/;���r��R�����D�S�:!kW@��_ɡZ^;�|��hP,&+{��	:��/��	]����ckhc�Qѽ�݁�F�.�b6�x��
q��ЯL�v1v{W�a���#���{���G �b�PV�B��]�"��A�|Ⱥ B񺾾>��⮇m��9HA@/�xi��:�L�S���ٞ/B.gl�\��[y��	�|�i�Or��7����	$ot꺝T���jd-�=��K�K��_�� 4������K�����8�h��cb������V ��"�zc��E?� �#��v�ǞͨY�UC�������W��3�/'���7T4�yx��S%���ϧ|��<�OY�'XM��J��4�,h�Eq�,ft��f��r��=E�9��82��Tb譧��M�EfT��y�z��Еc�Oݬ=v��6�rB�6�RCzZ�]k0����^��O����g�2����6`y�]��{N}��d�����I�e���76�&9��8M\<_Y��e�ș�G��70�*7��r�Y���^����;B�@2E�L�֥�G_8�)�!�u�� ����"��ȋ�ȳ�704d�le}q�p��}5��*��:��#-�U��dH���/׶x5#�m�j��ePvp�~�^������ʞ�?_�mT���FD_�Y q�=����.pv�νRǡ�k*���qh�@��7�)'� �N �ܪc҄K�Wb<J�Rxq˵�T��\uJ��\o�=Ie{��t��U��;LL�C�KK�3���;���z{��r7~�1
V	������f�쬶��M/��C��A��Ȼ;{K�y�fu�,�(����\m��x����=��24���n�W��O��L����!���ì�����BŦ�MH�� ��aŌb��|A$X�c��AD�O�J��_�7����H6��ɣ\M����Ư���-w�g��	�J��������QqqqD�Eč3:���)" �/�KcD���ئݍBO���q��yHө�dp�����c�;�|��n�y�#'��*��<Dp�2�-2�KI����b���?�^,b� �
[ow�����Z��[g����R��Ȍ�����ʢNJ����^�j�\��[Zc`�L�_]��zY`ǘ�t�p����_g��_�z����'��r!�_�{
u�LdV��7�1&�����S�S
�������������ӯ~���y$�0A��Δt4�rl1mlQ7!��co�]ZZ�f�����Zހ�^� B
�l<ѽ̭�a�P���k?
�z��ʇރd��NN�;���mY�FCą(s��exc�����h~qQ[�ˤ[�Mn�T����g栕Uυ���o���ud�($�vk l����:�N��J@Qe��.]�|99=]W$����|���DS��Qc�hzr�D�]��hO6F��	O>�U���P&�l����8�"��⁰�0���m�,�|;���/�Z�hި,���&�ȴ���I�'@�p���>:�=�#�C? G�I7�c%aWc��)V奒v
�3ҤLI�s��}K����o�d�e��3pyW"�.�Ąy��Ӟ^^���N���8�uKM��y��������7>~��MćJ D���]���f��2�kRf!�^���� 7Mز�oda�o��P������31}Ɔc#"G��ƞ���T&9��Li�A��]l��1rk�s��j$�␬tp�2t��-�r�-e�yόx]������^F��2�PE���.��k������|ۧ����~��!{){<5N�b���^"��k��m���c��U�*�b���P���Q�-p��e�n)����K]R"��6z�7�~�k�h�`c���2���Ә���̫xh.�Ю�����%F���ݲA(1�e4���wǴĥKYfb�%%%��f� 8��(.�+�V\�~ְi5�E��-M�p���z��r7T�0����q�32�w�,,��A�>�k"�팩���'8=5E��K�SwvG�t�ŮG�.�Wpx1ܯ�lV����"UN�Cr�����;Z�)~�����Tn���f
�~:�pϦ��>�@�x�"���8��A�'��,s�������_��-^��-������ew�'�O��=J�el��/�a�(g�;��7]%����1޸Rw]��E���&2��E޵¶
	=�1X�R����������e�C��#x+G��k>3�$9m� {�����ON�T[������~�S�tjj*�O������/�>l�b���|)��^sQE��Ǹ �ݑ���vz��!�[:�bb8T��������[�I!����r<�WUIzz{��.d�(��I��c�^�1��ֳɟ
�<y��qc�Tp]���Znq���1z ���O�Aؑ%DО J"�nl�w2��DӄF��@��w-Y�!*������[90��{s\Z�͆��� C���*�;=/)�D������E�5P��=h��q q�ҋ�"���~t��!�D���M)�x /doo�V�@�.r< �Y�W���!^����5����e��_�Z�O��w������{��t�ݛ�v�-�!J��!1a�����ўW��A���� gY��J�Wm\_�}�8�����`uӕ�e��l��r��j��L��.h�Z��D��f��v��t�q�6�G�*��D���؆w�l���C��/�k�.�~hȤ��"=���O�&�iԛ6���x#>�����+T����y��D��ŷ��Y&�<А��^�l������^����U��cR��|Qi���0U��� ��wd!*�Ǿp .�����:Q�L ��M�g�oVZ.,�d
�P?%m5��K�3�y����0�qؙ�V�9r�3����0�JgQ_^^~�~�X����is��n:��N��R6�PP�g	�/��Y��MNN�]_�8K�+(B�E�h���7���x����*�2m�sxe�����!��$w��mn|�uϘ�M(�;�D,W'�� �@zY[��_�wN���@�9��z�Ys��EDp�))����Q �� �Lh.�]%��.�q�
�=SPÔj�C�����}��BPCׯzC����ʰ�:�S�P�� �M4�G	���W�a� 镍��|zS�6����%E/^���˻��LMyO7�m==tTF=�&��ާ{�ӂ���^F5|�c�����4Q�.���tQQ�d��a���π��|`��ge@���t5��O��ry�;p ^D�Z �����v��6@6��2ǡ�n�:�2H$ve���uPI0���
{�1ީ �Ey�;��񩈨����T!C�Y�+)u �j���X:O��1��0�}Y�H��V[�����n��E�ʟ�t�U6�4����
s'�o~yYW����8�xc���##==nD�)ej��Y� O����@u������[��;J���Y���s�������%�&o��ء~Wf��}c<ژV��ck;���`�(D/��잞{@��׹$5��N���-r�L~��D^��f^?�i�i�A��)\=��!�]��n��qv��w `���!�sXl����s���lK�Y�Ԉv(��
{�O� �oiъ�^z�Jx�[�#�|P3o���jD�S���bccc�蛪]�s5��!�����A�4���S�yvpyY����!�ur���|t���IA����<ѐ�m�����F�����B�J�?(%��H�ಗa>�)�*��}4bz%�F`���q��rt$�27��v/).^�tn��@n��~��n���NkG ���n��?T�5+^A6QW��x���g��y�ƀs�ZG�Z�w�� ���q#;B�s���4r���� �e6�[
x�����X��M�P!����;��ixZ��7/��)^�O�vk��z^�Y��������/ ���1�+�V~D������C��ɹ�S\����c��tG�����s��/H>`aq�X``೨��7�7��w-A�q��V������ ����%�j�4���d� ����ghNQ镴.����J��8Hu�aN�� -|��@o�]�%�!JJ�ƒ/d#6�q��/��wou�^�Tx�lS����=��R'����� ���s�	H��#LL�u�l�	�'Bx�,Z3��<��f��v����I$��A�S�	1Kߡ�%��@��k؇��E�1Л{���sb|�L��� �A�o*jk?���| �ťT�c�ةO�Ү/w�L�q(ѫ{�iy���nO %�OI�� 7Ź��c��!���&Y�L[@��*�;a�tl�N��A�ɞ#���r����)�V4'�<Z�p!B)����K�f���F{''b��\�
��-/��PP��(4P�m/i�)P�P.���Ǌ󤧹SҐ5��mT�:�b��\��~I[D��~8��,���,��F3PL�%���.EX%�coŋ���W:q��0E�T#���S
4{��/䵪׼=��9(���$A
I�UO!��J�i8xx|\,<��t�(@��b���C�"����&O���}��50$3J�,op����@���ֵ�Ѧ&�<��2ẉ�Z����t�13`t�W�Hũ�����Cddd
������\�)�|9�9����1h������^���� �9�PX�xɋ*����v��vU�p�36�ܰ`��nKHHȩ�[�	t�P��K� 7�!}6~��ThEI�n޼��cz�~pFt�V���nB�h����_���(Ͻ�<IR~��8(�|����f`�������i:D�wo���䲒sq%����\ƞ��sAc���i������\D|��{���8�K�ƞ���\;����Ob|?-����i���҇]o�x�>l=��az[�B��.���xs_?ߝ�}G�e�[��Q|��w�+���w@�ކ��)���	��0�\G9�'mK9��|����~�	p0
p1�䨼�z^=�*���ɐ��K�L�Jq'�o�\�)T:Z0�F�3������Ŗ}�X����-5��=e� HUw�`��͛)MMʴ|�(�?G�~UN���D+�I��aB�<iD�8G����2 *hOEI�400�O1��Ki�L���Z-R�S_�~G�5(T��rrr�W� ��w��%̨U�`���]�.���l��˴���g���jM��g��Ѧ�����_���R+`��K�y'n���O6��4�E�X�:��x��ld`Z�!!!��Â�G.+(ht��f9S�U�d:R��������yy�v(	u��:Ͼhn��՜k�+!�QP�,Z��O&�[�>⤣�$|}�o���m0�������b�i@�-��j|�e���T��0������$��/������g~;~o	Zq����c�}JqG_<���Հް�٘&0�V�8�bu�W��G�z������V��@|ow�߀J��uB����:)���?c&���mnn��I�(#�J��ٿ���ټ�ѧ��ӓ���pd��U��S:�3f3��C��n���L��MBB❶�|_\)�Х�h�(���6�����(yo�q�	N���h�.R�&B�t�͟��?6�;{�l2 <ކ�v�@����S��WF#����JE�m�V3	�4�x69�=1a��fϕ�kL풀񯮮�V[>L����Py�2�\��:���L��{��j���V��W��o1�T����~�t��yb=����,JS:�	���M��K
�G>���?Z�`5P�s��t���i��۩���?�x��B��%T�W[���g3-h��3ʚ(e�?���ld����#��ņW�^�sE7��D��'���G�����vZ^��I�1d�8	%�Rb�B�e����2~o9���`c�&�z�R�ġ��bZG� h�{�H���g�&#�ֱ2��i|@�pf�j˶���a��]�i>r%ee�Ui��&���-��^Z��2�-�~aZ�l�c*%ݵ6Y�XU5�.XڀKv(�� �,��@h���3E
i�t�����������?���@ ��(r�g�_k@���;9�,��ө�<f�=��03�i���􅬍|��5ȣx�y�6J����G[?m�|7�l��$p�LV�Ł�)�aXxNǱ�R�4�.3Te�Sq}Z���~���Zx�,�-8�^�~�P�gRISmIG#�+/S0B��hD�̶����9� �Z��m����G�ITە־[]j��Q���{�׮��v���ԕ�ѻ�$'4b�7
W�Ҽ��$gLU܏w��\�a'�ߏ"HHJ��8#^�[b4�V��-6���Q޻�ߌ����*ǡ�H�y�;U�e��o���q4�n������ݘt�"	�yT���C�S��\��}���l�}��{t���ͅm��i=Gtw8�y��=ȴ+�Rc>��J�����x���#�wrv9�s����gU14y �ѥ���Bj��oı���Jǵ���<��� ���9w�<i��D�
'Caaa��������v��r��.���T`�ƕ73�y��i	u���o������C#,Nk�k]xg&�_�p��y:����bQR�e,�R�#R#�91��4!?w�r�|Cãq5���9uuuh�W}�^����?�����Յ/H@��F���E���uA_Hw�bc�nς�f���gH���0��/�[%ԁ�D��TM׉�HA�=%�n��`���`>*)3����e�HN�����������
x*��2w(��Rc-?Z�h ���S�黾zU�0��11F(�7!�o��)�Nd��fޅ��
���w@��,/ȣ���&ct@�m>	9���"q��h�2��_�:�	v��+Wtz�.vv���f����<�H���RM��898���J\�}[��⌡�˷�a�u� ���V� �ҩS-bo}�� �u�.s�֌�+6e|N�`��ÄW��fbZ�Fa߽r&�������b�7t��������aȵL�Y�L>����ձg�}����v�4	p'���EP���"�&S2�zG3#h{��W[J��lii����r�����}K�jM��  ��@�p�w��)�W���7lQ��v(@�4�U&��� YlG�0�����G�/7����
>o�v�Ci|e��zp���� M�r�<�z����P�����u�@���HM��v�=zSp�F�=|Í������ �@�p�T�U�_v�#A�om��ҏh_lT{?���z.g??�p�׍tٕ�:P�9 ��T��nad�U>q�C��Y�i�C������^_��m��Hˣ~a��1�=�Ҧ�B&.�Smn����oRS���3ihi#��L�*�ܡ{��������u�7�N* ���^��D/�����������֣����`(P�1�}��[�&������?z`��|��*�0���пvܤ���z��:���.%���.<gn��&�Mw.���c���z�5S�}/Χ�Ӕ�PFg�br�-Z666K�KKW��8����ϟ��o� բ�c�;`Jt�8�m/��M�>����cT0:%=}PM�񝞉��h�ʓ B
��[:48�4�!�$3��\ -j�4\yu�ݫ~0^�&��նP� ��Ÿ���~6SŧY=,w2,Y��<�6 LT%;�Z�B�R���Xy�1�=��dO����S�e���S�B=_��t@� ��Sox�X+�1@���VQ>nNQ��7��JUϧ�g�o�M�,_L��
_<��i��'�
ڈ�8>>~U�|��X\���f�����&�t�y�/6��}�c��\^� r�����{i����� ZЌ䥤��I����^KŦ�&�R=���{Z�_&���&d��� ���)�<�Ī���:w �d�Ps�s@��B�j[��I��!�	ך�*�'�����Qr+q���E�������X�Ƨ
PҠ�9M��_`7m�����y�7��MZ����K-�4#^GRu���LY�ٛ�f9ݐ�*+���xwٻ��(xK���+�:��\g���%��WvP�3�x����E�G�l����[��3� �1�k6�nᒎ�2u�tW]�2CV��+�������K��>p8��2o�C�C�95��Q�r�i\[���,���0���i��� ��C��\�1�l�9���K��ɨq��#-ҋC�cz���}AW&�����կ��&_��S�d���Ҽ�&�o���ή����6���Vɹe���[�U�{|��5��ds��v��L�e�s& S�zՀ 5����p�Cbz���&&������!JJ �O����~�q&���b����G��`�xs��!�� ��t7Wz��B��`�m<���~�$4f?�-���ɸz�N�+��K���j%��s��_��ݾTt�z���' ��EZ�,,�&l�A} ���_ s	O�1t����KR::;��O544�������Y ������ɩ��[4M���J����?@L����`l��#LH�����Ƽ|i��Yq�Óϙ���Y��$�0�+����v"���ƆL�$+�\9�S���؝)J����� O�V���J5�Q��׼�O?�C���SDw����-���*,.V���8Ӫ�_;��k{9�����vQ��N^8��� R
�O�UW�+k�鳌���?rRҖ0�9���`"�FGU;J�M�t�GLR�#Wkԕ��l��������X�y/�.����%A���[
/�,��-���+2v�j*l=҉P���14��ɩ5���{X>(ܿ���KkF9� ����wr��
�r���ݏN�(9��tߙ�`��� �{/lXe;כæ��������>mCCL�)pQ#�!��
Ͷ���:�B�o}��W��r�c�F}���ק�]��_��wtp��4Y����t��ͪ��Z�U��UVV^�b?�D�Nk+?iF���&�x'�ȑNk��㘪+���  �@��:��O[�i?(%_����ǲ]_�r:�J�ȼ9M؊��=8*�!@3�s?����nY��|g�&�JLVU�Fj�(��L�n>�B��d�X�����c��ԑ-5���� ^���[[�,оx�$��&���i䱦�b��. �wYm*������ ^�z@>�M��1)l�f�쾂p�
z�����?�۸�B�E�4$7`&���j|G�k��L)����A�gg����;�w{�$����rr�&7//�6���س�4�o'�mf@&<8��H��CgI��0/B;�.�>�'w��q�>�cXc�|~���?�T	��n������'K��(W�ِ��g�On^͈�rn���C{�`~�=ei.�rZ�C3�@O��`Y�h�#���Bx~ء��K
��웞g���)��4h��T��*�@Z(d5�������������Nȕ"�^������ni��>����j� �\�o�(��i"��7>�z����-?ڵPOY�Ӥ���� R-)9��,��cm���]�����i�hj膢"����#%�fɂ@�m[w���уX-�]��K�n�v�iT�OaKspd��+?���l(D9���ч���{�
򝾐d�Ԡ�X��;%N���q=]�2���w>5zv�������O�
���1�'~c��靉��;5΄(��h��'�����{�)u��� IZ�t�ֳ/�*1z1����_���s�%�A�GW9a��]���"�����X��о��"%4���c����Ug
�d�F�X8��ٳl�l�? _�	\�'���¶T&����M2jj2��^�Ue��S��]m����y��wX,�*V8�`q��6\����\@��+�q�s����Yޢ��?]LH;����醫�]z80�w�E�Y����1/�?&���?���¼�ؼc�"~�oO�{��Ͱ'�SSS���z��
~�ѷ"�ۃ���ll�L�ʧX�'[#;�i���́m���2�tG�/�WSy"Z����I'LՒ��]��I2e��[KE�rV�p�0SQu��d���sl��1QQv�C�Ug����z�= À�&C��ؿ�HVm<8B�@��6p��ޅ<{���y a�� �����Su\Q�Y��C��\�J��s�&u[A<
^�m��2���5������V+_D���8p�OeQ11X�.�ح�l����L������)==�Ψ���{�@$X�l�5b_: 4�ᶓ *|�N���p'!�.��Mz�OB����k�x���DQ|��\�fI�R RZ~��Y��Z���Z�l�ߘ��-�!�D[ ��L<��Km����S3��w���Rƾ*�!.�����?���F��m#��d��H���"}��,� � ���c;����v�oSn����������X��'�(��A����]�o"��?��y��ΜZ����m{g�_���^���C� (ȸ�rF�OF�b�u�����w�����ӏ=6փ��l�8��!u�7���o��4�&Vt]]H{�6%���焉�e�����g�΅����3���^�H�W�H�uj��|�<dj�!R������s�L[c �Z�,�b�X�#�ZUŵ}��R.p1���'�m��u�3��w�uI���iۏ,�g�P7e���[��z;q�ٺ�C��(�1�pzH1*å�w3MHx�s��	D�`YWA�y���ӎ�d�$�����zw�bTt����P��4t=�dp��%�l�.�DaΨ��jﮩ~0���f
�!�BBR���H�[��o-�(�o%Aqy���m��+��O�w�H�������fL��zL���20>�o��|��/Y`��|�P��0�����Z��f��{?aj!��۷��AL:n�	��4a\͌ �l�����Ù�9_�_&�O4Tч��(��q!�P�������\0>{(�������d���9)(�88/���#��'�9�%BB;E�Hh�Ǵ�:�q_0��{���nw=Oq �4���a�	�(������wҟ?.�!~v�w�|���9�]��Ib|~��:T������U�(5���3r뒞b�v�HBE�ty�^h��e��v>%^p_~��}��T�TU���C��ͥ���TWY>UMy��&�.~� B��)-��w��_B��[}��w�J� SqE��YZC=�B�J�R���*�^�� �@�y~i�f``  ��'N�|��ܽ6Ut)��ʧ�=1A����:D�k��v�>�7�hO+LD��E�|6�cpg8;=?����x�>���?t9lK�O"��6��}z#{𶔂B	�l#����Kޞ�v��� K��Ъ �ot���r´��ў���-���/�3g�m�zz�FG3?��I����������.Kоw��-\������%4��yk��\9#�uf��MP���[+eu6;����d"����Yh?����
��Ҕ7o�o�Y�'�2�&P����b�ofr�����g�ܴ��M�K'�.%Yd��B������}&�98X��m(D��B�۽�w��ʉ#�K��h�9�cP��E��%��'���w�/����y��'0���\�%ȝ;z`��ʇOq�b9&�e8����&���Ie������u�T�ZX�]���~>P��߇�� �����4�Ml��t�srptǝS-t���
hzs;��UFSUԛq��#��obl��t��7\��A7�%��1�a���='_�sv7�53r��Fi�P8�B �c�9�uu!���Sw�Hus���m�m�3�X�$c�
~���[u$dg�����q��˹ߊ�z_����S�ůƕ��b�k����A��V���,:`Z� ��GO�C'��>��V����
��M �;TU]�����Ӎ9΋,��7�I�n9~|� ڠ�騫�qm�-�'�*�����e�?��*��uC�JC�@�Ll7��(�9
`����ō��~=��(4�F>����:��Z3��HeM�cX�D˥�=��ڎ�@����?���8ύ�y(�.�R�5
&7>��j����z@e)&9p����� `\aE�b�i˄L`�6�ٳ��
�����:Ҙ?\���v ���Et$8��Kg݌�~<��"����6kQ���c�Å�bWVW���Us��)++�t�F�R3�r�������Ri�d@�@�[���E���q�w�#�4�p�r�D����!G]p �ju������c�ys~�fV����/@q��eb�ImR��.�Z�I�Xx�����D�Ϲ�c�{	P1�W2Bg'�m����l`p0���CI� KBX��KDb����n\0�
����!���&>]�5w�ǘ�
�g^tc��7��K�˲�EJ��b*�S���3���iw^�y�ҸO��g�Bش�!��d�3�Zr<�%׿��#����#u�߾s�@,����O������#�`�-Y(��ɱ�� t�~�n�ف������ 3��rޣ����i:��ՏGʁ	6�R/Q�	AVz�E�qoO��G���bޝqZ�90Wy{x��LEmFo�1q���;`LI�C��0Ţ�E��J�P:n�Sȁ�zo��O�7�b�:z�9@4n��+��E�8�Ή���쒐�)�����W;��l�B{��$��=:�L��J��Ó��l*  n'"���<S\��d���.l�n�#QOh6�c:�@UR�	G��>��3@�	���94�2�A�yǽq�o�_���2c<}M}I��d���T���5�Ǖ$�	|��r��cWii+��:�t��+��b�l��R��'����s��\�t�j'����os��M쌕�"+��^G�gώ3e����=#�\��z�(�/~tEDR	i:�[�i�$��Ar$%��C@��F��a�����|��<�y��c0��'�^{���.�+�n6,��H�&<`���ef���%�g8���e���·���U��VVy��9��٫Y�ж�$$nBi߿k ]:��i>ٟz��I������ǒ����&���"���t�_���������B�;��6��iأy�q�(��/V��N��L���`���6��2�wq%�f[���b8PVM�ke�>��qf�(#ro֛���8-�av �=���{M����Z>������AL��r����b��$b����!�΢���[��P�^6�I��0H��Q����j�eG±�:�>3?�,��3�;����h����[���D��/]�Z��Um���O�j�':�f8����߮�lo��͗x�*A�F>�Cm�BW\��p{������ P�������k�NcK1R����@�kHX��~A�9����=��� ������2�n����C�͘gG��_�˫����(�P'^�h���T��m�C�
0�8���%�Z�B[A�!"�=�D���B�x"@P�q̖����J:ٺx츂��B����X#tycV^&F�䠬֍�!�S�;��GYYY��� �ҷ�2����*'-���2I����>:4c+`�L�	AvN���i7��_�k֧�9u?�_������l��Y��W�vy��8��QOOOB�e����0�ttt��ɗ<8�o�LLȞ��
X�1Ǫ���8<~��ߥ���'t�b�z����z��� �}P����u�24��2�!� `�v�̽�<wRQ9v�7\Qp7��?Q	���R�Ӝ��'�!))�5U|��Ho��4��@cr��:�-c|
t�ҐG$]ݟ�H.�?)ᷮp�;!S���=*nmƅ�}]i�x����Ŕ��w+����%��n:P��G�ˍM��c߾E��F��Ӫ�d���r�ZҺ�Z�Z����	�U�����C�ŁT�@�%XH�/ޮ��;�M�r���y���
aT�:}�W�а�"��ma�I�2?\]�,,, !BA�P���Ȁ�	P�@�IH&�A��n"ns���F�A�I�x�ӵ1(p�9��i���W�uq�OWm��9V��!��Rjv���r��)@U�x�,@(���\�mp�8�����@����oܳ�?<�fq�@ �K�2v��'�N+��^�\Q��*oK&�Vne��ayeY\�����go���|^ʈ��y��N�-�d��Y�\诲�[��.���M��?����и�q$�v��#?I�db��c(;zF/%�gWQA�z
���L���{g�ūW����ݞ�k[[�Rd���9��ʫ�)V��~Z����;:3�������Ά�����O4�����n�"�+�m����u2���W�*�m�O�	������L4���;�[��|f�-4��p�2�صc�j�ʪ��wPG�,�ƀ�4	�C���} o�Y���^r�����L_Fu�{����.=O_?c�U���n���K{Ճv��Z��X�4�_R���U���d%�wQ��_?���s�D�QZ�3.�"��No��OΜ�<��|21S�L��Z�_/�ܝP6��XH�`ך*F�����i^�
B�A�,=�����7>&�vZ�V��*�^��h�PL�-�bmN�M���?���DEE���{�c���T���[�e]�IQ�J�zx@�1gxX�1��[�,�OAR��uA�+�,�h0�L��h�S�Q��<�Qr*�W�F�w8��<#�R?�8]�zR!�����[�)�� ��[s���v���8��qQ���O��N��#�i�ݻ��Je�����߽3�@�JP8W�!�[��M8N/:<<LP) ������L���&x���^=��^���M�̿��$"2Yu��Ą�Y��?��}z�Ҁ�l���������zӝ1��UW�H�z0���$���l���/�=Ugo��Q����ý��|֗'҂�יVq�Eݟ�3�-6���PG����1�~��Ղ$����w���mRv2���]!��)ᇐ�P��*
�!"R�ק|�uNbb������b 	��V��t�v��=�qLW����Cer�jQ��			QO�
8))�T�i�5��ڕԶ[`U��9)e���mL�@/,|8��C�n;B�B�QN��2],��Y莁�09�)AMGW`���f'��i�,{{�	�F���ޜ�Z$Hm���z;�b������J�=!�p����DHd�'�j���Ƶ�H��.�{��Z@�c�'r�ʁk�Z��: V��҂כn]t��;v�p����}��iɣ�N=r�O��_/@����S��'W1-���E	��C�e�9�dw���cE�ڀ#ϓ��ӲʃW��������d=���J���|�攼&�^�M߬A��Ȉ־�
1�B�UTp= �2Q�Se���ٍ�:�G&��+C��:*�?l`��V�Nqsuz�Ҳ�����D�o��ma\E���*��8Pr�e�	���ee�E��MMM_����A��<��QE������zӋ� �!~ʗ�[��!��RP-@�
�]�"�ݩ��V��).�����}���
$Su��;+5���y�pO�S�W/�tcj���Q%����nEe�ʏ���r'���ԣ���>��S�^o�^!��o<?s�y��f�>��?�O�PQF�L��������I�Pхnո.��}���B����F	�>Y��	��' o|߷��}{�!��٢���3n��������.;Ŝ�OԜ>/��h��Ԕ��߳�O3����y�ECb'�,��6��K����a`����ʶ5�4�nX2�su���O�\�����즋�/��9���־�l��_��݀��f���v���3#{t�ՍK��	�t�̇ք�_3�RT�'@:�F8�e�Yߖ)l�XR����V�vHVx�zS���O{�0�o� ��L�U��,hSB!z���qe��I*���:}�Y�����D����3�!�\�w��^:w���y��!�oʕ����><�Ndqe���T����Y�ʐx'�<lg�Y8�y{YӺ�~�rm��LW�Z���[�c;}D�K]2w@���"�ݫ��qA�y~�	�"ɖ5X?����B���7#�˫[�c��}�:�ThKw"yV|��&lޝ����痛P˗Zy�j�\��X��/�S?Zr[�m����8Pkk���B��T�^���ꂧ�v�~��EI&�o܍�N��K��6�
M�<T/l�������b������r��I�z2}���߽�����J-�X���ez��@��j�" �
eîk��uEÇQ�II��֯G��ĉ5�8&
�ٜ�D�o_=��s��2rSް��bu[���@�O�e(h&ȜӒ�5���Vh_D���<�=�΁U##G�ʊ�%I�����	=�b�o�7|��[��J��¹;�}��Fq�5X;���O�Uu�}>g���|��ŭS`T�`ޑ��y45�cJ�-`�C	ؓ�$��:�"���^@M�z�� )?�Ѣ7���P�-5%�����~�_�� U�y���_z��ﵜ.�PeHeJ�����A�iO^x�e��'�����]8ɶI%�,+������p,�:a�H�>nJ�zF*CC[�����k��c^h����j�'�l�f[s���u,���:�&�P�5C6w�O&�z}[x�[��?78�\����}"sOU�:�)_�8k��#�`�>�u��3ޢ��V�̃;��y{��{Uhܸ�a�a�9�I��q"\���<WP��0��w����U�U)E�S��Ӂ�����ޥ�-:X6��8��CH�c{�N?�,��:��YTG
tb}F�7d���I�Dc�9l�0�F���yx���."�;6ړ矿�j,1H���������m�H�H
m@H�i@�B��ʚp��.iC�(�,I���M/���qGVx�KdZ����W�����9@���]���+f)���U�,���DB�\�!o�Q��{�wa����t�E�"�-�<$i��1�+Tq:��]hKJURc綜V��ֈԚ�&7�G������Kx��mI'�~/	N�F+Ey��䒙���2��m��j|�����W1��
Ub�bQ4���s-Yw/��k�, Iae�r
tG�Ǝ:�I�@�h�ԛ�~�x�Y�j} 8���2��WTĕ����w�6�H��W�
�����i���['�yA�,��D��ϖFK��j~�&���Qﾫ�_�7666��׳:Yk�Gf�H��/��w�s��I���	�z/%�50�+�b����{MNy��"A��6  C���QH�i+z��a�.�b=A�Y]�Y^su@h.���BW���P=�c�Q	�N\:�Z!Fb��:v�
�1E9a~�\5�y%8����9�G7h�g�?�jb�^P�d�����Hu��5��Eِ���_�v���$�.��"Zh���gUKt��xF�j���-<+/-u?�m��^��{h�j�Ĕ��kӚ�&Z&[SB�wvv��{�����i#�5����]hߘ�>�G)��܉pz�iQ���*��%������'�
x��Ej���B�g}0tM{�ص���Z��D�]}���">h4�^YY�qq�y��L��ǣ>�89�v//����P������j�o�22
���� � HH\JB����d�����i5S4��(!���sr�*5X���7.#���/j�q�YNA�]���U�v��E�[5EyK�����)�1U74��bd��D|ŵ1���]���iճr�UPئY�[\0Xj(����%��b4m�mS���_�mm�V����YD�e��&�U�H^�- q�����yq9���J���?`�]N2e��=��u�hҼ�JA���]P����M��;>4��:� �<�M�.~rr�����4j�Zu&�ۤQ���{��h�NG�t0t �:��ODc�dC��6Q@���]/�z�����-�8�������nW���g���YKC8˘�އ��dw��� ��sN���I�g%Z5D:K䑉QF�$�e/�Ñ���W.����OA��VTac���K���g,?��9�n�^�W&�(X��KYt?��Am/�}Q11B'<�1��]p���~�T�m�t��k���$H2�^��D0�r��}��~}{��&laڤ��f�*���������Pn�xb����V�^��\[ul��qQw�����Z���뾻�"n=����Ľ?`���I���j�]er��^�Cs�eR�T�0��h����]Y�6� , ���'Y��yB�.�@���
�u��o�3���؇4�,��L���wQ=;��S2�;*�!ɭ�D�NQ�?9���(�ڪST�(��g�#õ�v�:5z{�>�t5#W�[��f}X
P�@��Bqk[[Nks ֫���q����`��1����,Ho߿�0�Dv��[�@1��b��Iܨ4�6��t���&/�\���z���K^���٩�<
��8oV�x���R��]��u�W�b[3�]aQ6��1���M{�XI	�}Ļ6�� ;����\�.&�Gj���<���@Dt\eeL�Ie��p���8-����V��A�H�,�Ȱ������=��>v�(9TRR��יn����A>�y�u����W�V
� ������6o�ԅ4Xr�٬$tb���y��Z0��t��i�����������زM��,���.�/��6�D���������|��Ne�2����B����*p%�ׄ����8O*svͦ�/HKl)�5w V���Bނ���uuM[��޽�P��+(�+�&��C[�����֞�t�Φ�����
,�E�ք�L�R>j�Z?�?>����:�������K�Z�P��J1جƅ́���m���M��3H�q����I�?���8WP�h�����C*�clzxɘ*��1��u���� ��XVV�7o���5��)�1��/��?K�x4ϖ���<��V����9� �~�Z���mv���|g4}���~"���u?_ߗ�^��K2< �J�T���d⿂6�그�^�
�!�i��

Ớ���ͭB� m!h��~}�.�u"��yt��%�B�Nx\����&@M�O.]�cf�l��	!(h�� !%�k�C�$�XAɺ�y�9'Y�TM�_.�5�7iHf���f=-a�Z_޽?׌�\���W�kH!.TF�F�1�F�j�(:p�m��xuZ���q������
�����2��%���I�WP� \�v|�C�M����3.���		9���|%V��)�*B@@^h��M�m~^�G�<�Y������[,��C0�+@n"��MY�$�Ϭ��G�9�����s�L�F=_uޥu/.yP��-�����z>:��!$z]�ׅj�^ > K�%�>�F��
��S�|��kɃ��M���ad��K/1�:�âDu�n�on�0F{���F��&%K�^i��a�J�Ir� ,����l�S���(Z�|z�IiO���$�F[��p-*Y^~P��m7{~^���f)��X�����oNr���Ub�N�YJ�V���l(�����]8$3Į�� � bݽ��f���񡦥�7�RLQ멱h��{�
�.�qP���l[�ˀ���_�Hޏ����{,0�X6(G=�Ŵ���l�ymLTcv�6��,��˙���y�`�º��u ��Y��S��iZN..�Z:Z`�D3
+**^�[^y)�?a�Z9�	��������`%��$�6}	�)��h�M92-����^��ʴ��4�d_%f�>�Ara�е�#w~�F�	��B�
��v1;l��rH���1�s�^0��D��+�-��F��8�J��h�ài�~�����.��#��ad�~�Q6��O��:��4�Ǥ�k�]� ��>�;S�֓#Vih��9t t��A3�vl�ׅܥ$xx~���9��(ǝ��O�M��I����IfUn�R�� �Ϊ���(r�#��H��v����d{PP�2���M�}��0�~�@c���,9���R�;��	�}"�!��2mS�|���_�'�&�sn��^g0�Q�i���h���e�}*tA��N�u�`ܟ�^Z��7c�S��va/W��T	Ph ��,��v�0ښ	��F)��eb�J�~|_/�e5�.v�{Jd�u:Ql<�"��i�RZ:t��Aɣ�%��\�02�B%�BJllp|:��@=���67�V(���k=\+�&��r�a���$�k���#�G7N� �#%%rZ@�٫1/I>>W��G�ߛ)�\���6X,�ڙ��g��,Y�EMC�����%���.���c�KK�o�}�z�y	���	���a!���T�B^����M��D�m�eNj*�0N��c*q�k�	Mxy�U&�^]����@�T�se��K(�1���1�x���T�7h=1Ԕ��=�Y*��+&[;������v��%" ��h��l I�F=�C`t���D!�]�!�����}������K/��L��b��� � �eJ����ވ�@u��w���-~����l)��&a`�6��i$�ͻ����,ߗ��r��RA�I.Ԙb��eZ���Gm�4�L���
z�0�� -�j� �
wQ�ʶÇ�W���#�[�݉���Z���4��7�qֶ�����8�\�b]m���i����@%eݝ��(�UF��A5fm����Oݍ�ٽu���-�l.�hj+-���\a���ѫ��}(^Zj�'������A�b��?	u�)�s�d����6Pe��g����Iq�"¯_�m��<=� ����:����x���CΈ��V�����(�m�P���&F���*4U ��Ҿ��TUUE��v�hd��CݍXU���
�f�I�8�����M���4ť*���Y�܄\��B:Y@���G�� ?s���L�?�X��RHhi�@ĕ���TyF\�/��Z�I� �Qf���7���47��t77#��~΁�>�~b���D�������Ww��"��!��ʉ���Nʾ~%�*n�{>�0;��C� ����YZaA.����8��E~=/�����GFF�Jzaf,�h[�נ݆W�MG@'�+�R6޺i��Ky�6v%ͩG"5���_��!��z�l�ڽ'���a��q34s��o�������qT�P���TFM�����M7V����W��׼,-uǎ<h�ݳ�=�(P�Z����eB���$\�7`m)K��tO-��`�Od��X��$
�] :�W�-n��c�c��ݫ�,RS0��F(B�qtl�GN�.Du��LB^S)q��`.+%3)���c�hT��P������ge�|��J��L RԚ�EKlS��3tSSSs����U�5.AA�C9���0;>��bԥ.�E��!�S3T�%2z�D��;=��<Ř������܏v��3��H}\x3"֤��m�n�n����7�J�_]�����0��d��c�s2������,�F�PK�8���2)����?���Y�3�萳t�L�f�"Ham1�P��7,�ۥ6ܺQ7���9mR�����bS�a�����-�ȟ�#���Hº���N�WOrKQ��w�: �j�ųȯ�{��<��Mש����״&.�5z�l��K�׏���Q�H��G)��)��f�d&_����\]�[�t�X+���R��Ȓ��2�_Q���PC�ǚ�F����{;nz��G�J�Ê���u�_�4AU*1iyq�a�@��Ta�`����`r�sx���A��R[���T��tvz��x�%Њ��v���9��!"�F���8���>��&���}���h÷n��iO��P<����A�����@"��!ƴ��>;QȒ;�%�/���;g{�ݸH�!Rw�>J�N�<�FPsN���*|�H������(�L�M���	υS��.� 9�,ҽ%5��ͥ�i���)(0�YE���ݻ����]�Nk�*�L������FW����Pd��b�-V	��bsxD�0�~N#�)e��i/�jI���P��^I!#;����8wsn�fgg3}��_A9��N-��S�l��u������	P� į���������4�  �PK�&��jU]M-y��.���ܨ�T��]��3w��ͱ�&eCcJ^��������^A�Iu�al���!���� S�N��s �Rr�'9���hպ�u�v�r�n���Oܴ��[��¸ğ�@	�<��q&�҃��e)�k����(t���y_�]W�t^���{�n�r��U-.斜��6ض�z�d<N����e+�."]]�U��Ҁ��ZyEP���Fxz1ꨋ�9C��5'/A:�`�gr$��^m;�k���Rlw����*d�ЦA3�u^?�ym�o6L+��:�*���;�6�clq�֯_<�I$~d
�C5k�.1���$ �5\"��X���Jz�	�JJz���'A����:G/	;Uy�<h��Xp*����x���z]�sYu���]r����	�,Dq�^6�9���0���u�4�w��*X_>O9�&|L$/� ���Qh]r��bm���\E���|0v)_[[{t�/~�v������w��������K�*�DgM��M[�Dt������Xþ��Љ��3�7FM�SS����ᦏ���\}ɫ�D�sۛ����4ৈ�s^��6jp&����o�5�4���)u��X]2H���(��0�����i�����w|)j�.�@ˣ�z^V�Z@�[�s٩"o��<�_/ ���3���wJ�}��{���p����[NT	�c�
�g� �>�֟�����޷�dR�!9��غ�9\.��1��)|,I)���c ߁���h�I�`�|��<����n�,"Wi���}�q�Ag�X�0&��O����RG)���졹������ɶj�5�����әp+�_V�@B�m�&I��'a.T�ot���'�������(^ �k>|x�5��ȯ_��΀��Z�6�����*��T�%;?*wu;?6�5X����+�公*�.�w/�NMM������PGQ:���K)�n�w�o��D��@�<Z]��8GÅn�4����{���u^�@<�$k��xDLY��H�ˤ�W��76.HII)��D��)t�Lm+(00ӱq��z�Cc��#����▨{�)v��>�IQ�XG�O� �W w���za=]����l���� `B�,XNN�ፍ3�+�^[�mm����� 5���4��q]���V��;L�|(l)�Z�$C��=tyR�c虂��Uxn?~♜ @@ñ��]�&x�R��>Z�\�����Gu��WK��k��s�G��OM=���ݱH賴��}Ʋ$��y�w�T�1�K}_1:9p��2ь�R�G|��ܾ>��z��f9�G���,�׮]��#{2�!���+,\٬$�����bbzO�����f��ʄ���o�j��Z]��)]�c��y��*���[��5u�⫚���&2iJJJj���� jH)���)�Cx��t�A}J|�S�ĨB�5�*�&�.�,ӞR�i��M)-�<;�6Ԁ�p��� w�N�#�yR�a��v(�P�L��`/Lgڼ�����т�6�b=tNY��߫/��^�kx��;i���^C���.�����O�'|)��54����� Gq���X�0��T�� ^(,�F�w�:���[60>�����Z�#��L�Lt|~~>~�b��:t恺٩+q����oz:��	֝N�9{�U;�)@~cO�k"��5P(�@�tSp9W�	�E$tU̢��������R;Urguh���w��=.�� �~H�N���RF��*�L���V����=#����\1/�m`��	��{X��Z�'�M�3gM�bm7�*�+�x�F_w����{����J�����#�=M�Xr�s�R]�b���烙MY���Dt�p��E����c3N�
� h��I���-�^���&�ĩ��V�INd��-�Ւ�L���p�;!!����B<ِc\%+]�X�!T�F�d�����/]ʶ�G�N�>�Ú�*c&��#(Gs������ǧ�v--31l��L<ij��A&�Œpk��uВ����aR��5A5�2��ؐ��2l�!� �VX/�@VVV ����H,Ɉ7�w��_�y�e�4h'mnp:���KHT!��3��ط0ڢ E�sv���[gS�~�@���n��~t��*�=zM�����	"Ү�A�!�����E�ZZ���("
j�?��
|n�|u���&���U�c��+ Km�`�_5�����L�~(���+J�vo9��oY�O�4W�.IP��T�0�ң�d[|����P�V���`Ogܤ�aoб�J���4�. L�	��E���}UFB}�7�C,_R�yg�w�����anWyE���sss���RA���K� %���Kt44GF�'O6^��*:H
������7��\ �<�$�3�#�ohtTg ������T���`����d�;�7<�_p�k�*��Y���<��
'�u d�	�<�8�U���C�o��;8��nw`V��͌P`�B�{��7�P|P�ӵ�(W����m�>kR���<����]�&:�p�( ��Q2´�o޼%B�zy��!��H���湭"��ḏu��;��F�PSv~�66��z�Ӌ������(L���{��G'�Jq:u|½�Wo��mV�\)��O�����upp��z蜴UԵ�kdd���ll@(P\�k�R� a���p�}�JP�~��|P�k�fTL��mU�LV Y�,�&GӞ���c	<5C�i�g7��@'�|]Ԋ���J�"��h{e��h{��_��c-�3@pLR����~�_��5�"��B"�`}k�>�/m�r�W/BA�����u�X���2wƛ�2�7�B='�c��4�>��������f��������bu��D�䉛�k�"����RR�w������}ܔ��
nm������w���4�y�뷿�OH���}�
��(�0-�!^�Ͼ��,rt�qe  L���:��T�ϓt���Y�����W�s�	����O�-nu��YW��㗉�'�Uno�k��BS+�ٱ�������n�H�C�Mhr�s�)aD�$����	:{�y�T����ח����r��H����jWWW�C��^$/TI�]dR�V�0^���ݔA��.�C.�^��#�����(�����OO���R�Z7�Xv� 햟��j�FFP�Hʬ�tQx���������B�ί��<��0�#'��N�����R���A�<a��ˈ_� ����̌z�R��ޟ�����m����_��ʭ\ֺ�IK���[[rY��;�����w+�]h	��0�sm/�_$t�:IOCÞ�Ӗ��֐݃F�4`�D���9�xm'8'��t:�����u�R���,�ǉ0(?��ŏѵ&�#5���ם�����yM?ҫ4��?i��S��UUU�DDD$������qݾ|����S\X�S��E���	4hƜww轹	��N����˘4�s�=[y9晿.Z�UR���YI~C'��D���IY�����z�<�W{]�Q}���.3�'��#P��R��X���>��[pY���kh���&W[Z�q��?�Pow�}��f��H���u�89��ۘ'��c��Qr��С��sH�)��X@o;<S堼:>ɒ��x���N�#�O�X#%.�vrr�4}�[J�Iy&]SS#��Ύ4��p���]c;<rT������-&�ئ@��H��:�s੮9^c��)ո�,��к+A�MrvVN	��杒A���ec�r\��A��0Iӫ16�4�`���K|8]��o��X�5�V��RG)�=��	����4:1�oqu��G�� c"55��C��O�%�~�Ee�<4����J�����g�w�	JLk&~d���Dia��@�F:L�I<��6D{|�r+�N��+[̕�:��@A�y(��xz�ǵ��ǯ`0l�J:���ccV�sdR�<��|��#��of��_xh��&�1�Q>�k5!	�U\��〓P��N�v����-=����3�E�Q5�?k$X_�Ծ{�f�&�-P#�����ӎ;rT�z�� S��f��:Q���}��?�����y o'z����]bbbi�,
%�"qWB@@��t������q��ڵ?���]�����t�z�f^���o�7u~�#�![-pX�����>��0[Vb�鈨����|�6I^�g}ZF����^3�X�'%���%?���@;�Z&��%%�<�y"V��!���F -�-���'�#Y&���q�t5�=_֠��̌��k�tb�ٌF�r��K�p���8��Fbq�kpڲkc�KO2��n�����;��1WR^�b�s����s~~~�,4Q��6�k�@%�IB9�Gջ����e��:�΃ާ�&HO.���
ї��,�O�Qq}�Q�磞��n���k�o�v-�Wb�4���鎂���5c��Ҭf���Sw3 ڮ�9 �	�r8���+J�t����������?���51����<.��T�hc�25��w����rp*kR(� _��	�L�;R3�k�ɫ�u��g��22U߳���*)�L �����a+F��~Cߦ�\c�D�~�5CC�?j�!5'�>��@背�{�Ne������_�:�;����jIQQQJ۞!�^�1�`P����?yʡ�!��C���ˤ�66f(�������'���75�A���Rj���k��>ibk
���%�3SO�:���X�dni�	���K�=@�n4ʃ8���M��}ZM��t�}[)�Qک���:��"�V�S (��q&x�h����<�Ǳa�u�\������m��lQ ��}�!e�*�+�5U�$�Ӳeee�5d�IE��RW_J��1��F�`�y�_p؊U�o���T�o�I��S �-���� MM�>-�%��gQ&
^7  �6 N�Q�m�l���?���hdoFS��la����|m�&(����h�\$�'\!O~
��gąν_�<\kG�4�f˲ǣ8A�cc��~�G�\��֊YF���7�Ʉw4��΋���?���w+��r��;��=RXmI��ygP���n�PJ�uyttoM�/��[��Nw��z͸:<:.3�@�f'�� ,���\��?g��0݂�Knok� 0 ��(���D��(/�Bל""��G�0|o�S&�L��n H�x��6�]�]�D��K��O6��/	���d�bT���j�~���B�&�`dIP7�yID^������8��B"��)��|!�!�6�Z���E�����	?�y�ڹ����殮��3bOZ�x%�O'�܄�4dW����8��N�MMM&ו��2�,7�����׍��/�O�6�!�?{�U�Ӎ����13���������Q���D���PJ��:4jbi���N:�9��w�9��$Y5n$�{ʱ2�r @�4����g�zmx�[r���iA��y��fb+�
��)��[�Qr����c�o�j_Ix�ɐ�� ��t)���ߘ�� ���q�k���
X&b�V(�q<(xUQ��H+\�����\{Й�;+�󕦤����,���]��}�|иA~���
9���dJv��lbb�����j>5����d�mP����󌗉�|M%8�9[5U��������M�O�c��P������mh��  ����w��TѺ�������7�/���3Õdߩ)�X3��\K������+���S�h�g�H�������}v�=�:,���i�{Ӣ=��VewR����E�'�V����P��t��t�r�Ó�!��c�۝A�e����#S�- ���쉃z��kSR��īL��# &�a�&�I=����G��$�1YA�U��X�Z1	�R��y��JN��[���p�-�C�����Q
S濉w�D�٦�{.�C��o�q��P3Oyߴ�|����L�uF4����ޕdB�9:���b�8����"�%۵�����03{*?�vm�@�ę���2^s��D���p�LBs{�qZ�Գ��񍍍����[��|o�/�lw��M�5]_q���O�U�cjr]V�F_�x��2�SL���oZЛ9`�<$�BE�^�z�y��ʄ7�F�Z�'U�S\�*l���9�J��R�s��6ڒ0�����c�F"n=�"��;2����_��i$ҡl���k�-<���tAP����R���Iܽ
C?F"�9����A���snnn�?,b��%܀I��1N?@
���@z��E"d��ii���LPt��{��3V��>㓚�\��Y<��^�U q����.0�:���$��	���r�|�ݹZS8
�P�3c���_���Ȥc/{xxԮ��Uk��r����py6����U~�@2���]�ƌz�W:(,��TO6��sۻ�T�a��>�z�y< ULl���*�3��0\ɢ�����-��@"`�-�y`cRkp�1�Y�4la[ZeÜ�IhS���'_ښ�R�+t� h�S!n���#',f��߸�MGn��>Z�YY��k	�t(rd�q~]��A;\�=\�_��<�%��-`��KD��)s�Y}���8F������������;���?xˍ�O���j�C�R"����R߼�:�H���`��w�}�p�X��%�s�m~�h �h[U(aǳ���V�U8���L	?��$^��C�[�a�J�V�'*�~�͓��0b3��&Cr�m�ڐ=T#St?� v�^����#�0)YY�*D��ڀ=�?go7ra�Їԅ/p�����ek�ExH2hMڸ}���{�Y���R�d3o���OC�sG\>o8ס�Tt���6@)#
�j��"x:�pd�t�Y����V�L�J�!�O��}�Mf2m,��U�%:�II�8�7m��Њ
������[{{��=CjU�Ȃ��e>��t��j�y�{������_ԢG�5yZ��жR��IIA@dTR�7 &;�9�Y�1�� �¸�o炤��������)�s�M_)�B��M�p_#2rq$����ȗ�f�_%�b���#�����dq����s�!�B�_A���&���-_v���;J����s�
��r�?��6E��?nA�|xf��U$5+���$��Z����W�o�B	��[,<b��ҙ#F_u��"dX�F�Lu�&L�UiSE�-���хF���V�li����7r���_4���B� N�����z��A�����W��a8u�-4�3��30M{ذQ%�b�J��p�"H1?0��9��r\��k-x��	S�yo��=E�}��_X���Mq�A�ia�ez��%+�/a.%m�W���({���0�[ܤnf���w�I�W����I�����f  v6�e��o-�I�S�g����^H�HBw�j�?)v�l޼G����$DN��7�}�p��K囬����sk��u�H�"�| ��?�|���U�PD"�ޤxi�ono��$a���N��E�	������C7�Xqi�.��0���>A3��y���B��_MNR?�WV=���{�F}�N���9�~"�+@���<}Dw�iz����܇
�9���>ZT�ԓ�8`I�~�d�8ڨ?���I��MMq��#X6�R��K�3+<(W�I<�a���#��o�!a��X�Jbŗ��h�ݚ�3�֨��6j��TZ�ӡ`v��eE�_I��N(��"yA@��*�}��G�h��~��E���D4"
`��m�FN�C�Fׂb��ֶs��ε��ʞ�.J^`WN���9M�+�eC�j޽< տ]"�i�:->Z�r�끪�����d��vs���5"""1�u1��ML{����.��K�c9M�Щ�EG��Jы��P=65��z��AAo�ϥ�D.����w�R�q�# �C��]�����V«o`���;�(�8w�
~b��K6�$(�%.ҧ�n8�,r�y�F����b�)oVX]�e��wO9��J[_K�|�U�u����Y8;0/E�X0�I� '���X���������V�g;_�^"!����c����E��[�~~��֡�m��M㘦���tY�|z?9P,ֱ�tK�="2��K�0Ƞ���U=��1+�9^9�w)q����p!�����VhP���%�B�r�Ҡ���P�vT{ �P"/����o^���R�l�ɮ��:[������t�Ö�'(ׯuE([C��'�Sь±��*���Fq���X�ߝV�P����N���\I���MJ�G�݋MIs�q�L�Z�+Ѫ�Y���?��Ȅ�]D,"��M��[����Ƞ��� ����Ѷ���#��:�s������z�?V!�����FA�(l��u"]�z]���id�:��BC�\~/7�J|V-Њ�1+��p���������Ty����|��Ifb����4����X� � ����Ŝis����`Ͻ�-N�T�\V��l���~�lH��b�$5�����B�0~�L��+x���>��|�	hc����ٿ�0�����?L]w �o�?H�"e�
e���������u�Z$��"��ޛ�	�{�co�w?F������<�}_���>�纟�y�������B N ��0?�2A��:�A[j2I)E��c��!	y�䅬OJ�r݅�9+#eA����x�bI�[�ۇZE��V]\L�����!y��ȱ����/�0Cq�n��ϿZa��sS�V���i� ��(�����D�Z���T�I2H������J���ӊԩ�7�XZEj�O�N���%9�"�i(>�Y�>�&}w�Vc��c���ʫ����G��lm=qq)I=����F�J�X�?�7
�Zpl�U�����8?�U_�{W��'�D� ��.�h�4�A��[rW�v�"�<��R�55池��ۂ9��`z76uy������pb��Q�?������f=ͥ�t��Fp2U�E�������ra�ΠW5�z�����cV���W���"n��%I�A�G��-�N۾���%���|��g���ĒB���\���u�P��l.�Vc$=�
�3�� 2尨H��d�u���Vdi�w��9^�!����p�nYW��g�a�c�E��E����N�o�y���>6����aOq�Q�U���S�p�����R�K�&Z���K�N��rw��ݛ�6�/��ι�}@�r wKd�SU�����	�ˡs�{s�%���V����\����}��⢓0�mq�� �;��4bill�3*�%��/�];]d̹�z��_�6��;h���ϱF�����kV��:l��:�^b���1�'m��INX��3;>��}���'���N�f,(�P�������ߠ��|���oJ���k��e#N�.�����#�����>p�����F�)���:Ar���:�B7QL���g���)@%���N*~�����#f�����Z�&���Z�����S!EMi_���V:��#��Ag�*��l�*m�Qz:��Rݲ��?ǀ��Q�>��KE;��ay�S����_�����W��R��iR�}�?2�o,)��xa��Q~�������+z���,��	��U����f_<ߝ��J]��+X�.i���BEĤi��<�d�ykng�;�2��ZGV8A?ft���p/5��oo��ǲ�U'������s��q�n%�wwu�v�׌C�)��wZ�1��H��E1Sc˿L���"G�1,.,����mF�?�{Z\X0�X3��9\�p�W7a�Լ@/Ƕ��M'��.�|ys<��<F:�>sx�$���0��W��l�1��|Q��#���0�$m����u�X�ګ�)K���-���M�>�Yl��"�����m49{9�^�s��-�r�t��s���R�o_<ӊ��D���a�G����Z��>��S�����$��%a�����K�
4�Y ��~���hG���=� �Dٳ=�'����7n܉e�*-5�{c��I1���|����)ނw��5u�Eh�-/{u���� 3��{��9�H]/��Hmm����Oyo|0�ߤx/u|�rxq���UQX�h@c��������[m�:�_TI�>����l���H�s9V��0J��vN��J��3��O�U�Dd�]�u>��c� �Cq��b�{y�����+R@�8�oY�`&�٫� <��b ;�:�U���=�'�k�}��`ɱF�PS/2/�ݺ�<�����aX:���Q��vdU��z��p�CܡG�ŝ?sx��㎖��Mu�Ń�� ���(����z+7_����(��v5[[�����3��K�Ci���1�_XAO�R�������j�^�[��8�!i#h�*��A͒:[�����������\�e�ɷ�̈́�u��|�߽#�d=Y~��Q��q�m�퍌 :d�����&�ci��lb7�U��V�A���%l�$�-�����q����z|���:6��y�<�H�'C���m�l��=d�ª�D�c��KQ�����4r,m��	Y�@�t"+���h�2�����.�0:����~~8-�^�`�Q7�'z�_srڱ.>h�#X��"m�q�;ֲ~K�Z��t�,� �ǹ&2,�����\=�U����L���i����R�.����ݴs,�2��K�lw�˕ɽwܫK�71�&����n�O��$��	��)?�*�L4��HU�a@�P�Ő�8�u����?�}o���[���I4FA��
���z���d�uCܼ���H,�hr_#�����m��bF�o֓}i+7��st0�;��kk%&׳�C��х��J׊� #��S�{�[�=�RI:)����ʊ��5�FS�\�e����q縀�{`���>�Y��U��vS���){izs�,[��~����Um.o���~>;�T[���۷ɉ��w��ߗIWN,�����h��9�Gb���O�E]x翕�(݉H6K��'w�wF�k�����.E�|�0t޳?���>v:�'�f��?0j��o��7��f�z>�=ꖧ bk<09����AN�x|�&,���Nd����'�����<��K���-�4��)�	�W�g��'آ���쿲/�͞O����c���\J��9��B�Ky_1����H�����������:��@� �l�<Z���P�@��qA�`T��"���Ԍ�dVUv����P��Uzn�9�UzN��ÿ��\E�0�v9��D.�,
����Ӡֻx�w|ܠpHG<1]���8l�35s���x��������h2�O6e3�خW�p��'|�{��tll�k��B�w�7���[3�w:K�u,p��|������>TV&�;�����:w��j��Zwi�)�*x�X�\x~8L+E֐���MP
֜����ݫ�\=<�������?��A~���@o}}�F�G��(���D���
R�\���9�+֞p�+i�T!C��I�N�<U-]ɫxM�+������i	6y����Z�N���:��G���_�:¥W.�V����:Q{��1�@%w��%ӾC��o�|[x�0U�p��]�P#���l�bDDD[�ws��X�\*�*P���FFFzg��
�j�x�zOq�b/8|]������t�.�CK�b�VI<�&��0�G���<0_�T��έOn}�����B���V��3��EΔ/x�b����bxr����ҿ�<�ĒȮ������Ci��l�˰'w�B)�GG��]��������[�3w��wv�k�R��'�lj �yf�K��dp=�W
~n��ZhYCS�*E2�j��C��M7Й�M|]ǀ��WB\�7"J���}�)�]VJ�ӣo�xq@�G�d��`}�����N���I���iV`�ul�K�r�޶׺ �j�vi��o�ָ�o���2^|����[ZE��������3���Z���� ��0��r�"��LR�<�	�^u��ષpj�-Y���lfث�� �9��ڎ��`��>�ۮ��ԶuU��^�����$��:9�U�>t��ڏVn��%���Q^w��#��!.�(��z���	%�(f��ş�v�g6�P��x%T��v���kZX�}+�P��M�NP��M[b���'�(Ӿ%*�ϿJDd��ibec��]#���Tg8���n~�=�v\���x�{@�W����
��o A�3�(�_��g�ݫ�B���LbJd|�-��vt��距�<��xb]~|����e�����\���TogѦ3��Ȇ�x�Ig����dC��ً����姃�>�6��Jk2��� H�և?��9��.o��]C���"�鿭؄x��*�7\i�w^R��AG+�p>U!��̱������D�!���X^�P���._�?�2��V�-x�%2;��5}������ݓ��5���b�E+�E���hb�Ϛ^NKKВ���f\0}��6�g��2:��2)_ZMu�5�� �)�QG(A�ŧ�(k��P��H
���o)�*�Q'�����U?���������|�׆v����CX-�
<ݎ�^��3{S<:�R��ȳW]s�U�u�5U�^���=���ݜJ��3$q{ 7�*�,,�ο���&�7����<��Yu[��gG��2\��~�vU����Y��ӻ_ϳ����(������+%�G�[����e�fj�\�{i�+�E����{��wm�����~jjj3=��pq3�_E^����M�G�>ۢ` jW���U��Z�sasw� �u�lP��B���	�RW�;��΀����`�:	�����M�3�X)R��%�	$�Q}4�e�_�-�*ɫ��,f��w?���ԋ99�^�.���b�	`�Kߦ�B�Q?ֽOI�u�ڿT5s#|���}�{�O��G	`�v�: ���;y&ѶU�xcF����vwJj�]+t�� � l��v��hy���Q M�<j���*
q�]��F�Ѹ�,���=���WVV�:�˟���Dp�ͥZm�8P��5>ma����>3�A���#S�����^��h��D-��2�<0�C�^a��C�{�JF��`P��X�M�:)�&!�D��pM�q��_kk�Q̰˕�!K��˜��m�x|t@��'��(�$^�ځu��ۇ��Ź-1�����1U+�$�!�����6lP��g�l.�=vY��}�k2ds�=�حX�J�{��L�ׇ%>�
��>�BoSnpͶ���)1"���YT��<$J#�z��bуy��px�s�j`1Dm(U3.��rP�"��ݔ�nj#G�aI���e���/�c���z&C��C_҆
�-uL@ُ��\{K�~:|�C��-�X�N�S��˓�ޏm]V:�9l�=#OAI����+
���谪�����x��&�D\��ѭ,���V�a���C�Zk3 ���r���s�xǖ*XF%r&Dʎ��S��@r߇>�[���	<g|�]���r�A�QB�k&ѷ������WRM޽P�w��=��}w����>mGk#�k|�}��S:��؋u(�T���;���P�f	N
����orM]���Cx4وE�Wk�7l�1�yz��~��p5|i)�E�O\�CiX�OO������#�,#ܓm�U��I��A��,�? n�^+[Ά%�����,�����($1ٶqП ';{�z�(g4��,�Y���F���"mA�RHnF��񍍍2PB��+�xG-��㞈P�@�>L��P�:Q��I�7�_����W�,��s��ӍԶ>פ��'��<���iޑ��ɘr���lk�bֹ�f�9uy�kS�{���xMM_v{��ѝxt�kH�m�*�o�����p��?��2�lŐ��9���bKw�Wd�~Q�-r�x7{w[�n"�����\��vY��5{�Cȑ#�����~�_豰��1�h�@[�%����'�ƍ�^%���5T�Γ~��Y���E)�T�G��qJ����8�\)���'��d%<��dO�Z��ѡ�hh��������_���
?�8� �/M�&���23��*=ѻ|�~	�R	}~�άC�����{�6��p��s��U_��� ,�8��	 �,m�[XنN� C�xJ%�x�cϤC�xarR
8D��?��YZY4	���-�]�BYl-���k�$^<~:�M/�0�5�PDإ��e"t��s�Pz��S��&\��@���~�WYIC�̂�a�]eP3���?��{7�<Ѻ����). �>�#���+A65|ɜ�
L�[���7��Ɨ��3s�|�ʼ"Bl�X��:��Ӆ��,�A������������oҾ�UX15�H�"��uOO&���J󤨴�*3���و_U�Ề��� .����=�6�@-�Jш{�&��R��|ؔxД@ {�ǒg�#�9j3.���p;|IP���R�eS�+��p�4`���{�����0IC�V�N�D���H�>(�����iR*�9,��n����H8Ȓzp��n8��$��[�Y"�/^y?h��)�D����k$(7҇����$`�W=f�͎�k�x;���NΠ(t�3�Ƞ���;�8f�{3Q�������_�<��NW��zU1,w2C�f��������swM���~NX�?ܔ� �u���؎�\;Z]�f� Un9+;{L[�@P�"�P�m ��G�|ŗ�ķ��Fp2k�3]ݑ��-�ƂvqL�����n}6|�ݚ���~��IJ
��DӮMY��N��ϟF<7[��8 �j^m��:��n�ƌ�ݾ�bm�h&H�����W�b��d���1t5��
�u���._I�Y|4��A(vC"����ȥ.8�q|��[�HӐϾ26������Q��\��th�2^ޛ�>����W]{r�2�=u�Tv?'<��XJ4���`~�H`
�����<$�`�,�iJW�W���b��3*?D\ځ>{Se\1����� x��G �gq�'W}S8Kx�哙�4��&$q�����<��J���a@�cl �	0��8�������W zEQ��Hu*%x�fs����VJ8��r�9�;�S�,שO��7��o�#�4 �cO:{�^a!��r�KF�m1�?1�5y*|(0Z����9��n���.*��r�̠�A������:���qT	)�'�<����0K g+�s�p�|��3���`dPE����i�.���(١J�u�1	�:`jf�hQY�u %@�	�V�y��r���}� �m�B�abr�9���K���Wj�)�����*^b֢X���W�6U�,����
��"�=�T��m�!�<�KI� 5 ��98n]�)}T���d�W�2^�KxA�|ff��	d��X����bdz;��T�����k�~U��b83��F����V��)�]$#{"�QE�)�����h��'�\iDف�i�:@`�T]�u͇b�{�˰�������{{MLR�7#�A'���m`d$�,ыpw�EƵ�p��fO���o�%�&�� \�\E���s!��bO�3eX��0�*�p��s2A.|�|u����I�G+,�!:!��R���D�D�t���v�\ms��RG�Ē��б��`1��	�o�h��w��g��v�
?Nb���@~C�	>h�3��җ����K���v��=`%�F�@������/����NáYy���^`9:��WhC9�*W���~AL��'+\$ Ё�>Y�9=$��㸪7�e�JK��>\t�:�6�/��p�7!_������<����s@A�$
Wr ��Q]��)��I����u�.�����@�����s
�o���_Ck⁍�х����ʿĢ����vkpW�W����V�߈v�<[9���_/��U�K�5)�q%̊|�Q�{��R��ng�7 G�Ұ�ڟ`;����d|��ĹuH�umT�y�Eؙ";V~��(?�^p���[�����R<����%������'c��C��s�=�K��~K붠���&�TU��~�X)v2`>�T�Ar�6�Ü��>k�����Ү���]�ȓ1;L!W��yزǾtF�O���V$��5���	��Ȩ(J��J�1��Owܫ�={��:�\9������8�k�Ve��h�rG3s���N}������0�jm43�oT&�A��Bo���r�Z8���^۽=�U���G��߿}[*�.����8�ZR+��=�@5��x�z#� 	\����M���b����L٫H��oJ��Ûz������A_�J�R��0\��S9q���tzg1W�~��Suri�o!8�ψ	`2R�$.^��^3���XQ��Sݏ��69'�ݓvE�7f1��4�_ݪ1�xȯ���>pU�=IXa'Ш�z�0���5��`T� �^L���!ШDԫLp@nQKW���(����(��a]U�দV�v
�П�Ӏ�C�˟O��}��Jx@C/)T���Z�����Uw�Z��0��É�� �؃��[j�%�ԟ��l��&�¸ve[L�g�c�_�prq�c[�K&���989�B��j�@�����t	߅���}�~��1G�N@�g� �gz������[�h��!��x!VN|�m����ޔ�u��hPTgT=҄B>��Ʃ��8	AA�����&���w5�H2ivv�zH1���M���555U ���pm���9��W�������S1�	q�`��ga��l��,�uw��
8�@��d6dh�ki?[�h����f�9GM2g�SF#�^�r�}FF��Q���E�_\x454Ƣ	��A����Uq����,���H���쀸����I���,�z���Zw69nv���
�9DY�זA�3�ڟ���a|��X��Ӝ�@���?��S�Cz��|���4z�i�(<����WݍVe����p��Bn\:��m��p7�2L��Te��f.���5j��i�$�h�u�I�ߠ=�������9e�!ڼ���X
k�p"��쏬�W�I0ŨnL���hd�)�?����ax��юL����z��:nB����o<�l��Ms��j57�(�0ɒ^ʅG=f���R�]]]�S�p%P�*�W_��^c�h��<aUfUz���$�� ���<�W��|q��yN�eQPPD���:��YD�U@`��	� v)�8&�N�$E�h���~eZ#y�&�qos��{����2J�t�*}[�7���3O��,�]���g/�	e?彉��)G-Zǈn��
�Ņ���Wɬ��K ����qm�2Rͮk�����յ�r#�E�|1�!@{��@�U�$��ܱ�/�@Qr"�<���]+R��hx������
���Ӥ����4P�}N �4JNՎ���h����D���8q����l��Wн��剛��8�G�HIӕ�Ӟ�솲�CZ�~v�t�*^%҄��s�4���c3��l��K[�`����I�����afgLQ�ҍ����5l+p�����B%��V�4�V��F�4�q�6M�t�+��O�6Oy^Vu����H6Y�D��������9ˤt>�y���b�A�i����2��|ד��m�{��o��ȼ�F&-%�u�9���:y�����h�o�ø���G�$�[V�ҲR��!&�Sh�\P��Bֹ���pB��3m/?�b��j����v�T�t��E��Dt}��5�7��i��}'�y�J����G��p<�'�<����QL�i�cn#���������[��FF!L�	\�>snv"��=5J^�L���&-�.��d��	"BP\�J����X���={i�+�Gl���M��)x@��Fw\w�#��;�
�Ea��nޠ4�Mki[S;�����vGa��ۏ�.�N<W~��_��o�N��@
���,�Q�3أ[�{ȳ~�S/{m��K�b�A��r���N�)�-T���~��b���Ch^�;��;gyo\��祃�%�Q�#��'t����?�Ot���5��~�8b��,S>.���h�K���A�!�a�{��B�-����8�Q���-���K���u����a�vE*�9�8�69=T�YX�M��$���(�MT�K����⶚�/Q���k�ϒ3�Vmn�6L,����V ��G�}·|FtmZ��V�ڋ?����aS��l��3�ڟ���0����*_�_-�r������ae-{�@*�mj���َ;�6�`!�ޛ�w�9a�Z�
���5+��Kf����yh�~����x	�	�L�FI�l>tt�?u���#?�lv�>2@B5��X�d%������Ѕ/�4� ��ɺ�{��:�	dD�W����~�9l��Iz�\���RqS�݇%���Yc,?;<�G ~Ч�:7yU�?_: _b���cM�^���M�!}~�='4���9��o�U��3G�W�C��T$Da<G�˰�z�:E�<^䨬����K��'��#�.pE{$.%�m1	�6��K3x�i��{�$ܡ��)f�o����GzH0>���.��xm��p2f�"� %�ڑ��`�CI���w���˟�I{���1�J��aP�K��m�+LA���l�ڠ�:��}��Ԙ�����ɬ�V�7�r�d#_Q1�I��E���(~�91�AS�u���[����#L��A��-�%�f�������{�-,؜N+����[L�1v���O_���|/��W��.=�ڡ�#�m���@U���Fm�o�d�*��\�UV~�������،�j�n�?W�K����59E�/�6�tt�iQ�1���'��<��`-}���Kb#y&Y�k�b��oY|����#s�_�k�	iVI?u//�ne�4M�
h���SCp
�ĩ�Jl�0��j|'1� ��E��B����U��!��S�B$Z��&�v�w�a��i�.�Mpt�%M>�w��bW���Td �d#���Ϣ��mc�%�	$#G�go)��}��1hm����Ԟ������YvŽ�8M��6�RY�� ��9��&<WsK��d�Y8&|G��5脋���_�/���:Zr,�f�&���y|�$��1@�O��ɤ?	7�[v�i���]%��)�-=�})�U�_ޣ�on~�H%y�Q
��l���ʅ��&uM�����������wRq�bZM3�ts�����ł�[�(p�Kucec��O�+$fg,K.�)���,�b�7���Q��7��t*�ו�s.'��zj�9����s��|���_��r��h�G�E����=/���qN�P�*���!'��!KY=k.N�����>im�+������<q�̇��@7�O����b����@ ���-���FP��![Gk>2���G�+Qf���p;}����ڋ�z�_y\�37�e-��+/��A�)Ӣ�������~8��|�m�{@�츑���`��p��hEv����µ9�SP�6^ar��q�}t�C]^^�n���QLD��_W��^���:*ʬ��<'WO/.f�(�N���� ��ك˩�_��vFG?�2N���y~ �K��ؔV�7���x߶$W��b<W�����:Z�Z�ڔ�9����:�>���3- N�'�W�E�)@������*X -f,`*�����4I\1�%�F�*D�Z)޽+���/��7mJ�͙;��Ԯ����QߚHLk��2B�����jW-o���x���)ۆv|�9C�e"���D��[ 9��y�<r�>��y�FP���}~Ӛ�_���Y�M��/u�f"�ڮ��	�����"MR�����t�D�SS�! \���N���h<q���n8sd.��(��Q�M��g1)_���]��r��!�\�
�]h����h����+�usKK��!��������Q����v��ŭ�Y�b�L���@���%έ��v�X-_z	�ӥ����Zwnu3��+ �N_?*�2[��Bu\��Yo����(	;��B��q$@ hY���׻��(�5WY��`0ڱ�l���PD�x�v���N�{0�d,F����/����b5&���T�DFE�!a�)�"u�{��6�ux��!%2{vi�
i�����2E�t�Zo(w��j-����w��Ķ6�b�W��ԟ�60E64-�Tef��^���c-J'r�0�rz�� 슠 ����2�c��,�
ob��`����E�u��BXS�f(U⎏7��s�c�����Pfs`W�Oe��Z��	��FU؃��v˜*~bZ����'ح�j�f��&~�lP|�8��N��}:FϿ�ng4�I��#ڛ��b|��"������p�`Pl�̻��Am��H>En�����������+���4P�˻�TI�y����=����"���<���-����U�M�Jq�s���-΀��J!�(u��d��u65�;`�������b�
�j��Y�o+]ʮP���p!��R�ւ�_�E ��q��D�~��^�8I<`�{#5$7�LZ%�����Zڔ��/0s�OfUE�G]/H6B#�T�;��}��&�i��g�O#d����-�P��6����[��o@>�w����L�3����Z
�H�"UE3��yT1��q!;�����V�)�iKa� _�g[Bn�J*Ȳ�No�z�����i͇	N��uŌ�T0:��ίQ���}��e+��/ H_b00�y�µ᎖R!�����y�!i��ᜮ��]��&�f&��'|=�o;��[���v!Dd5 �ٖ̍����[�U���:6���"|�Y��W>�ׯ�9��u���---v��%`���|��6�y³:eXR��3���)����I�����z�R��'�	_ngy��S�"UȤ�<��1��g���R��Z�����l��Ͽ��I���^��C�Kbkn����\��1��G ��S�Vއ8�� �:��V�c�#H�F,��<�c�q;`+VY��_�ZĲ��n�SӏY��8����5%��9�E�Z|�͕�:\����/�׏G"
�`Bt�i�鍡o+�Ņ{�O��< �KC``����=�s�C�^��b�o��'��պU͉��?����lY��M�Wٝ��v7J7�"ϒ���y�q/4X���v�`�#Ho�Ǳ$���Q�D���4{r�Fʗ�S��%i�z(M���Nk����ё�����/FGA	%9H�� -��G J�+;='`�U�<�+���?Y��2`��x��}F��t��o�#�1�a��6X���2��}|�99�B���᪼�r�.�e�*7�ׂ,��n�՛�����Č���;Mz��Jk�h����_t"k�<�+�
�[�8��o�HWjƮ���֟�����_#��s��ksD� \SG�>��������e;��<��@�8��8�<#^�Q��M��G�V��I����ނ'��5������v�'{�����|�/�[Q�����������Yv�̞={@@�y�)HT�c�J�� )��L"��\���x�IM>��������6�o��o������L��:؎o�?�M�@�y�B�����d�cH��_Ǘq�����1_�pZ�
`���w�>���;J��7�Ҭ�2��������A�����S-|B�/yb[?�<m�U��Y��'�r��1��?{_���m��Ό�]��e�.��4�GSrx'���'�v�x%�mËN ���?~2�5�������X��y�!*�٣���b[M��ｿH$h�%�m~��?�J|���k��yNr	�Q�����>BS?�ÂǰG��T��g�~Z;(��A��:��B�c�V��uID��W��yp�yO���ڦ�4�1��W����խJ�抔?�	(E��L�g<sVP)�D��S�r;�ؾe�����g�5�Y�V�9�egGQ�>5z�Ay��HT�QW�j��<$�E���"5?=;p��ݔ�"��%���\J/�����_�h?Bs����
M�Xoſ4�ѝ�Ӝ��ڪ9J+����_�jg..砬�~gi����<O�����x�������X�\�
j6�V������,�K�9=�Y)ѽ���W .3���RV�s�41�w�1�0E�x�?������t�y`�h�t%{�������~��~P!o(������Y�ҜPR� ]������_I�X�q��Q@2'������?�2���R�P�}�c���NN�ْs8���ׯ.,������v�ќ7�N2��M?@�?���&H	�,��٠�*X.��U�	���		��\��&�����,��(�Z��m
��f��P�d��{avRC>}�劋��`�;�o��%@�@�=�v�=�_?��k����E31���%��/��J7Pm���5��2rY��|!H�����kU?=��u�gfLүa�\EC:́�d��*i7-�Q�_��=+j�Qj�*+�e�M����M��	�A��y�g�k��@�k��~ D�(K��KL'�EX�"�;#��QC+��q���c�J z��}���w|����. *��U�?�S+���m�� �a���� ��,��=�� i�έ75睮�C��[��/Q���LOO���h��:��b��	���c�� 5�g�5�5��g��]�淐G�)�gg>]f��e�)8��1�O��PnL��:�l���5<����]���l�G��=��pe�ha��~��<��`$
��F��c�6�?��@�#@��5�Qg^��B���7����9�Gp�q���߭#i*I��͜W��4K}�Ӭ�e�#jw�L�����s?
��$b�#bWڭ��l�l�����Ȣ��|$�r`�2ͿBЭʚ]J,�Y�zM3ѿ?ބ�D.�&��wi���h�.o�/v��+;ލ(�N���X��R�t՚�ݨS�Y紜�������E�[U]�>��(]zn������ Hy=����=�(��Km@�)~����B  ��M������hdd�TFz�� }o2
���w Nbn�T�2-���mC����;rHJ�����+%�	�2}��<i�`��C�t�7��\O������+���d;�?�N@��	%vӿ?�l A�i���^Te���wә}���^�{E��$q߳$<���A�'��n����� ����|kо�J>z�ݛ����V�$�A�҇�ӹ�:-k��<�� ����힍S�;o��7})M�J��5�v��'�k���4���' |Ŷ����wV���e����&J9�z:W���3|B!C��%W�����c~!��x����LD�8ڀ��H�B} y�Z�~S�L���T��� =-Aa{
|��M�ԕ���B���~�Y2�H��O�� ��4��a O��S�v+E�i!�����Oy�����{�����l��*%�K%�Hs2���;jÇ#z��3�5}9� =�S����Ԙq�wB��e6����b
�`�?�ޘO	m�3B�1�@�+��rr�W�;#1�8�:H	W%9V+֪]'�@�o�mЊ����e�� t�+���9�NɎt�ջ\29��v��#�r���3�vÚB�c�#(���>:����yU� �(�VVVY��(�S�D-�ۆ� ��G �e�;�(PQ�hS�f��K>P[ŕzaS���%]3�L�?�%�b3j`�X	G[���0�w #n{^�_B�s�� �x�aWJ��c6���.�C��v(�(+L�qx�h�đk%�v�|�
�A"�k8���ޱ�oV%ܔͳ�ې�Aw��(deg7B�\���ux
^����i&50-.@�쮌��JM�
'x�n�򾯡�|�v�,Y�6����3�Z2����:����FA��H@W�8i��a&u��^xjJ	4��ehV3R`��&�{V�فʞS�2�
e��E��%Y^̩�d[�-��%u�ē	�}}���&�t�y#p5������`=6E��$���x��	b�O���6�{�=��M<��ˏ�a���_���6��"��
�BB�'�j�*��i��cD��_T$��U��c&��`�*�Fo�7�Y��|3MN'Y��������P����prys�	�8��Խ�QP�ޯ�rs��yقz��oP����G�1��yݶ$����M�J��+~�������#1~�KS��/�98RC�6�;� �=w�TY|'���H8>-�]��v���RЈ��4�hQ�%���]�s7z�����cy�`b�i�p,]�pA����l�D�aVN2��`�M)�>n����;,ymF�\�,��10�@W1��zJ-q�)���ݙ�߬�h�Av4����Eԃ�o�!����SL�\��ls��UCο��l_^�~�l�8؆W�}���� T�y���u�)�`���6?<�)������ �ٻ=��3;�7@�����eu��Ln�'qOz�DC��+��+>w��E�,>���O�*L�{wz��P@�P<��"�&R[��q���uAB/�:!W���wc��6[�ڐ�XT���֌��$����/C�]�v���hhcA�G�)H)V)��kщ?$�"T�H�#�����3\>�+;�����^�-��7V{aTe*WL�n�ڃ^��_&ڲ���t�&� 9!�3W�zo
�����/��'yȘ�1�Ml_ll,?�����7�ӊ������i���f��~G�/���j��JC ��N�F���B7�c�E�E9^���O�JT*����n*��؜Au2���e֢aɏQ�^�jv�z.@��)@E���NUG�C�HgN��ʈ�3�3�}7�[����A�Y��{|��̍Y?~��W��	��}G �~�J֖���W�<U�4�8AR���� �/ ��Z��t�͈?֚c��K��2)��~N�r�pQQ��+�^^s��_�dK���6竏���iNֽP��ۆ!M�4�d�5�]t���B+b��������۫i/LHi��Q�{���ǡ$��U�Q�)��C��c��ߦ�b���G���9���㍔��-}2i���,��9�#�n�(cM�=�A�\bkq�	�[��)vu��b�=GB]�����>\3���'�Q�!��)k70'���(ȹtg��bpd�'�j���v�V�M��䅵;�rw7�g+"c}��N.�B^&�%L�\]IFKE��OL�um�Յ��4�H��?G�Z�c+�ut���[�*�u{�~sۚ����_���t&>���kj�#yS��>}.V�}�
��V�Ì�u�eA��V��e��'��|�/68$�^�R��d�oꯉ�}�iW�C�-w=�ܪd_c��kf	n��3w���VM�sz:�����-�X�W�Љ|_qMs��_?pU���	O�_����rGv�jQ��z�� Q��xu�k��5����W+��W��y��/ζ�Sgeee��*���|�J	���6]:����5ve���E���p/~����KGKK�]���@��3U�/_��
��|��Y��o=�ٝx�|n�p�R�ѧD��݃¶���	4�MW;l�col�!{@qqq�����JT�Z<]�ݟlv�J�4��0�ӊ&)%E�ű�h���x�X����S��x�l�/О�6�C�X;x\Kp��<�zE>���Cb!�m������ !��o	�M�:�'�~�����������M�>}
B�;B���OG��o�{��ӵ��d�˰}�O�z aF�豮��%I�k|���^H�����!d�!T�ԮE�g���z�����Ż$t��h��њ(!14<��s��"��R�Q%�ߝm2_��p��w�ށ���<�`No&w�����)|�wX�q����$b��߭�1k}i@���hvj�kË����X��yLVS�#��$��W��Т{jġ=��׏��K���@��,v�UC�jj"�/�H!G��!i)7g[���&�HK�Ĵ=<<���]�`	��Xt��G�T6����m1�;�z,���v!��%_���k�Y�Nݥ�T�����3-)l�d��B�VW�kdi�;99A����V�W= "i]t�|��g��
%⪼�� 'C�j����/�f��o�10��w��h
���J���3p+�����+�K�#"�R卺�Ɂ)O�[V��O
���TS�ᆃ���L|3�����2������Z`1#�(@�Qv�+�sg�N�u��ٺ�����UA$#��RU�ɾU��Ew�>��&��C�h&�
Ʒs�����Yd;]��˃�h#BJQQq�Mן��ُgyF�������n@=��w�\��ǩ����O7$�;/@�*R��9���c�M{�$� �&�vp@^�d��ONNf���ԟ����0=@�m/��$BSиM�딦*����n�@ۣ�k�r�t9�%95�ֿ�2�#�����x�~东�l�7iI~�ؑ����s��I�����ј�X���Q����f����˧�_D\l� ���?�'��RXTE4��R˕����Ȳ_FMM�=Z��?�gj4|�o`����$tKIl���H�م?qT SH�<W�	 ��URd@��e�Q80�]�{�R��Z�.��b��S���C��] 5e��������w�r*e988������*��E1�e@2
��
*�s�DE@� A�E$I�X�JQ� X( YA$�R	*I$IF����t�s��9��ޟs�{�j��&3�����1�Z�/�h�S����;ݥ�%iHt�����Ne��G W�!WD71[C�iU55 ���R�֦^��Y�{͌���{BL�;�|���x�n��76�
�u�x�]^r����M�m�/�'���]�-8h��|��(�7�	Pd��5��O��qAB}�O�C2J:�"5x��A��`pS���ն�����
p�}d��hN�l���ȕ�u�_���Uf���v�up��ŎBo��))���C���"P��G���a��P����N�ԕ�����]�/ $���Pf�~�Ǉ�jj�?vm�����{9)�������p�R��/���6
�±�h���|��p l[:�����(Yߨĳ�7��g�����ff�,��i�	�o�wE{M7�J1�����Vq��Jiizn���{_^\z��h���,�0��5�*�NF�����n*q�`�Y!�+����'J·<��yݽ{�|�5�gֹ@�� �h��.Nj��-:�iu	�4��ÇU*�K=P��7�XI�'J"��7:��7��q��@I@�b�#Q��b̞����,���o\ؘnF���a����; yV��ǡ��	�g^\%����?��m�����F�ۛ[���w�!��D�%���O4��C)+((׻��i@� NMj]�K[y�N0{X��Ā��l���6L����l$�h���!�jOq�B���_���a��ڐz����=�	�k	
�Apz<r)�Z�vOy{��������P\T!�̶�����}���7�RJ9tu.���Dy�6A���t�p�N���ӟ��:z����������uTJ�4��2Z�/�N��%]Ȉ�X/yɩ��?F�q�raP,� ��(����]^�}�nb�7k��i>?~�Bsf�ʡ�rʻ
�֬.��͓࡝��,vd���0(���֬a>�t�<	rQ}����b-Nr�Z��9u�9����6�B�t/�!���<��� `�{�#]����]D�L���Ij*�Tu��/��t�y�g�B%����M6�^���* �;��L�����]���ڔb� gjC����u�&�nnn+�K�ښ먯�펽�utt��g��d��6�z�< 8��}	�hW+�2_��Ն��������v��}K��|��`��"��u�LϷd�����S��8
�B�;_U+����P8oC��p�?MKK�g�tV��<���ƫȗ��s�:�Jr<a*����{l�եw��D{�in3_;F��%��mv��j+:-t藽��Oq�o�P���u�ߠT\IP�ם{Iq���~­�3�z��nQ.jβ1h�uR>��{�~���	h����?���x�p	ڬ��mg֧��(�(������4�Tܞp��՗�{��:�{LX�Lo��������EU�><�s|ݷ����/G;I�ػv2�y��U�꺪��0�X7��ʚ��� �~��.��z���
��S
"���N����/*���V��ԟ#�|}g =�v��[h��l�N��3_{����(�TVr�0J��%��� ���|7�>͑�m �bߟ=f	�-:bj�k&�	

B��:٥gN�����������ݭm����`�_܂P7\��AGL���]]t�z�g�9��	,��(��<v�~,��jӗ�"}[[�� 9��赆���~�a�K6C���kٚ�H���A��4Y)�I��j�N��N�B4!ޝ2LIL�<�bl�\�R�P�N�������l��.hWp����Y�Ke�.�ԉg'��W�Q�, G]]B�y %o���Q� 1�.�\�+S�v���P*�C,��1�� Ud��)�n��9�L�L�2�?!.�Ƨ����;k]��O��$m�&3
v�T�i� c�[|}pN�%�����ggg��:Z�[��<�n�"z�H$�^X��er`�K�=�+�9�S�X�����%)�	ӋS{�������zܑ��<�2�� ���#�op�411A�+�G�窕Q�L�ϡA��M���90oA�������؉��X�QgRUJ�[t��܏FQd�.&&��5�;@F�?����������~�3���!UO�J�Em���$�䬔�^�a��;���٢��0�$��yg���~TYϏ����wBѮ9ˇF�o߾y0
�G�����	��p	 K4������߫>����(�/vbA�5]m��p~MCd�ʕ�[v�n���ă�`9�;>A)I��^,p�������9)%�(��o\�ˆ��7(��-\|(6�ڡ���Hɗ��15i��@�b_�/�]�L��1ӓ�0��~~����T��h��"�P�������*�ċ��VS��N>�S�c��w�b�QJ�ph��@ݾ�0p[��&����̇�F����/�όw�?��#C@u�[��{'�e�bR�)�-a�"�O��?��z�}k�CCf�~<��,��FH4�Ywȝ�؁36 ��}ū����]��n�?݉���(q�/���N�}��sx�]�9�������KÝ�.�~��k� �]s� �Q�0��E"����)1qq��欗-ٙ�n}���<���~|��>=�rs~��Q�f��^m�366��ڢ�:Z4=h���ޟJ����ڲ-��	`,亮��h���;MaKs]��mTV�(�]UQ�:/�ܦZz�u�H��8 ������W�v�(!p�ݻw��س���nq�V���@E�{J���4��	7�^>�%(%F����-���o�������xqq1�f⿽����|Z"]���'R<v#$ ���a@��a�@��H�)���'�ԙ�~��;��Hî�~.��FI�
=eA��g���F{�I���������2I�\��⑰�nY�0��S����=K��!����;���_N�8���+f�]�ho�vA /?8]Hq��y�Y�'��6g�@�'�/t�)J��l�~S%�tDT$�l��$����˖��b;F \�[^�07�2����u��s��},&xk�N�?;?E��Ժp�iz� ė�ci���$�<��Z[�iU��]�v��O�갧��C~��"��b�ڊHii�֎��ٳ^��[Z�RAA�oOn�|��N)ccc� ��a���}_��,����֦����k�P���l}r	�D�_�h���S"���fH{*� +*)�(++���馶�:���S!��pG�J42�����ɨ�>����#��"'	@lA07�4z>�B���0���ͮ]?jʋ���?�M����S����h'��+>�_M5Y	O�sjjt��U��.dX��
EO���v*I�&�H-.{���n�0A�Pq�������ʵO6�d�n���.�X�Ag��r�4�N���|�ɴ6x�{�c��f#�Y����I�ZI����ж:��|�;���^D�oș���u��6&��7��GBhE��a��ND����Fl��c��X.��?��:��_x}��0��_vTJ/�B���?
�Wd��ty4'!9yH,/�Q__�;������1��8q��?	�E�rt۠��+�.���Ru!`�Ƒ��ne=�=۶m�\Z��k��]7��8K1Kq]�b�/�E�C?&��#)��)��W��	)��`�����{�4��0Q��![dِz��U��R�����A�)�.F�qU��܉f���6�Ag+DZ�h,:����VԺ8L6�����_�n
	-�G�쵒cx����\gz��/�b�dz�p���0�oW�&���!,�<�I�12�O�B=���I9�/���SYC��m����&`X��J�>ϥ�9��ո,�ڨ�Ol�(�Ӄ���{R��7����8��kmà��68r,���Q���i��\��{0�:��䯓�N�:��䯓�N�:����ѓ�{��6��ݺ4��5��ţ�����t��c���������U�?w����͜�k�^��
����y�ê���_��o�o�p��N�[��V�~�����Ͻ����E���_	�%�����KJJJ�Vɭ�����X����(����N����&��������c�S�Ɩ�TTjW��ڸ�������I�N��&�n11�S>�md�uq���V�'M�V�'"���4uf �֟�YU3�u��~�����=�𵙡y?��>Ӯ���8��a��$մ��.�W�B��<�]\0�7��QO5j��knnn�.��Mz�`�}���ƟW�)k�H���&¼:�/T�:�pqq�V�2��l��ѝQ�UkP\�~]����8��:���TƂet�X�O���ǻV'X��c�=���b�����Ɣ����ʿ��K�/����8b1Iq�2�i!����Aܽ����$''����E�s����p�]eSS�e�����):F������!y�W3��{z�'���Pp�E3�;Mn�֞�MV���jZ�FT��@�0��������K E˭�w�ۅ��K��E�+[w�ۺ��e�F��[�:�L���ެ���?J�_	�%��_	�%��_	�?!�q,��zX�veeҽ���xh�'Iifվ�ȴ�cV:�?��N��8>�ƭ����O���s�*��_l#�o~A�?����K�/����K��;�$�<�R���9B��<?��˺���{�2>*h�c�;q�С#��B�_����]�_'��u���_'����I��vJ��#�9}P�l��s�N�|�^���������C�ˊ:��;���x�./|Q�n���N�U+��>��5M�z��bk|q���d�5�|�r�!�耧�����3��e(<e����Q�M�چ�s�Tda����!�%�{�8�K�֜yk��a!KA6����y���{��pݓ�X�G��T�y�g��"��):���z�z,~�GXNz�^=>n��vk<~	�+������b�y�ؙ8�Pۜ�3d-?}�:\�c�J�=p_��$���&""�L�JL^8����JZ�����ԑT�_3��Sxn���n+��D�����%8��R�ނ���r�@�
8�"��󔽐�n�\B���k��QG�c��_-����t�*"2R>_8��y�8����l�D��3��r����)��Z@!��U�i����ИCX/��`]�\XT� �=nx�U�9�#Ұ���a�Ǯ�Os?Wk�2Mk����7�S�����Ĥ��`��8f���s5
�)������8�,��o�n�#�ʡ��)��A{��o��֒7����Hx�3 E��k�j�CDr���ԏx<]�����H:E���oOi|�P����j�t47:���* ZD�\��QL��'�s�G����}_0*T?��H�El�!�`���[G�絉��tqr:��Ĉ��rK7e١���Oc-X��߮��!;E�l� \�_@�*�~&��ؼ������y����������J1

W�j�&���1qV�&�Fq9s��YZ����! ���U���-�3����_NV��l� .��dl�	��C�����tOn��A�B�Cb���2����#�����(����1��j�����+zm�4�&��ﭳ����!�]+B�"��_JRO �+�ayO(x�I�qe�9��a� sH:8�ow���h�y���j���\Ľ����1q����p	8ڢtA�9�$g���Q��v����D��L	��$A�h9/b�Qe<R�_k��	���v��}mNN+�H>��#I�f�I��b�wY�an���'w�"]�����r����?���sZ��:ϓ#�c�CV`ĜP�EƲ�^sZ�c?��i/l1g@�2�@8�g�	1���r2�b�!/u�r���p�u;���l%XQG��V�`�O���
�Ӓp�_���H����(�M���<�7Hr!���T����ɍw��z�p�_�v��,��>���p�����]��Z��_�E��q�UQ���Q�d.�G.�R06[�& +ޮw���,h ļ�)f�M\�u�q�Ć7� 5����2�"�쟝���7������!��f���,���S|x18C.���^TP%�S��8���,�F���w�<r�>��n9��J�Һ�bǑ��U|�!RL/ɉ����?Kv�(��9gD�j#.����,��i69-������X:�����x�w�������3��d���Zةù��,��(�K�vb�
ƅ��Ew�B�w:)ƪ�S!��,�q~z/���[[li�
6��0�zF�e|�Yh��B�6X��	j_8�L/WUp��v��е
ӂ���R�/�a�C�� <����gh�'.Ml�_����cd�m׸�J���l.��Nx��{6��. !�q�0|^�7Y����_'�\����Ts N|j�;�g�*%b�F�r�Z�KG�
���:�����.�
fB�����뢀�O:)��B?��bH�:�zV�̂�ܿ�q2{aԃ�U����+t�[���L�UV۟���8ƿ�J�i(F������ �%��WYp��m����a\sz�Z���^h&_\0�OF�t�@{
��	V�lbG��N��r����&����>�[�8Ym����b�?�ܽ4^�oGvy� �P��, �w�A��B^~���귰������Vy��<[��A�8J�*QӜȃ�������&g�"Ռɇ�OY៑���wf��'��ħ��$��〒����C쾝�r��j�������	�V~Аm
뺩������L�h�`c~t��t�w�3�M��>��V��8��cϥ�J�&���"������s �L7`��r���9��BAz�����~���y_`�>���M�`�1�ǉ��=�g%ͼ�P/�%(y����6��6ui�+K? 8O��7.�h���D�ry�Q�M-�zvo�M�L�y?� �cIc�b7��Ә��;@o/,X��y���Xd�qb���6ֶÔ�O �<��<}��%�7�fi�-��`��ͅ)O7XؽUؠ��\A������`�����a���s�R=�%>⛯�'���|g��H�ЫM/4�K\���\��W�}�I��>9���֦�ʣ���6���w� ��љ����k,����*��p�aFP�M�g�x��6�]DPO|=� 4f�:ݦA��u3����#,8���&��Rk�!R�V����=b���rWS�sL���J����A$X��y)&��~��������O��`K��j&&�����;�S���F`����DԼ�6�q���r}p��+�{dd rY�0�j�J���αm�c���Im��l
���!�:�g��%�7N�����L|f�1��N��z�+`;���������TCқ�0�Zd跡z�k�q
y`���i�X}>I7䔥�o�'�kz�Đ;�pݥ��(h�5=,������G7��Ɔ�c��Y�ۗ|]Km�7�k임�@��#�+�u������áa�K����@�G���H��Øh�=M�!���U�]�e�O|m�N��#��q���:���]a�5�Bhk@�e��@T+{�eh@�)��;�h{��'HM�ml���h9*6�z����S&����!�#1	�v���
��	�ȸ@��a+	�w����i�҈�ݗ�m��'fx��>�A�YY������v⵨�*�w��0�D+�Zr	���6٢Q�C��M6!R6��d~d.N;Z���e��\�s�YμfW�qW
�\>�����.���� �?�u����,�CO�+��ǧ�!4nm��pn�5��n&��/�;P�΁l��p��d�h�6�"�J���W@�R}*oB�,ݔK(3�}`���{�bsV��c���(�}��'�[�Ÿ�}��OQόb��Ȳ�b��e���a�Ox����C�hހ=�	�&��.F�@C �a�=��xp����'ۇ�������δ�|��7�6���0Қ��d�>����)��Oq!��D��,��k�B���rH�z�6��F7QE���d�À�BP����o��.��pֱN/�G��<�H� sK,��F7C^P�	���A!-'�;�Z"��� ��l��Bl��]��˴R������e���K#r�5�̸�������3����i�Z%�.�ݼ�߄���(z�ly�~֟}OT9��.�ԯ��G�f�r�&�hhvS5q~��s��n�X����(��K;��B3"��VD-2���"6݊ޮ���Sn���� 0,a!���������\�M@��+]_>����0�?��u(I� '�%�e�6w6�;V&4�	��";�__��u�)���_i��P�j���|nf����n�g���^�h��.���t$`���7���A-XmgIo��|�`�Nm���Ǟ':j��]���_s���*+��Jn�Q_�t�K}V�{���<�)�+8<��f��@^��@�|6�ЬCF�r�]�
��j>��р��֢艭!1Ff]���Z�0�z�?�tJ.��;@.짉����O�]{kA��J:�g=�u�\���k@G6⊯_/i%%�+<���b�#�Sh�	��ݏ�����lA�3D����~�j���RP�VH�d�<�����I�%
L����w��}�n_n?ǂ�z���+��ep����Y�S��R-j�_ތ�� ����3g��W���SX�˚�C�B�*�4D�pV�8C��{�޽{�/M(r��Al�G�[�\��.>#]+$:u3�'.5h_�"5���Ėk��vC%:>�r��v�f���'�>C�B�nW1ҙ��E<�����mL��pt����%0��)Ȯ��_M�q,Ԕ�a߲/�{i`�V]~�~����ǘR�A�p�3eB�8hܤ V��1�
C�1��ZI��WZX�>�'!i�*�<�C$����cx��#�YO _�;Ԫ/��� �Mk��{���@�n9r�0	�?��Ğ:��n�S�2�5���KƅqN���N��f#r�gwȸ��l6������!.�g��2������ܰb�*8����E���2{˛mV����{��Q��6���O�f�;�3̗��D�|�l�������N�ޕс"�	մ��$��Su�������(�W�7�o|�}(�3X��Dmt�Nb�q'-J�+΋�͞�U�����2*?�9�,q!�"�i��J)=y�-�Wi�?�ITWX�6r/a��.:���k��
Gq��k�r�uM��?�B������y0�����@�-IP��W*�}*�ȹ��!o�/��{�¯�X�����M� �S��
u����"���R,�R��0�]��;6���2���5Z��jy�g��e�ol���n��ij�� 1\�N��CF�o��>#�֣���,d<Q��	�IN�Ѷ ��~[x�6��yiݯ���rd��ŵ`x�]����*�����؆&�"��:����,��9� ~�G��������S�T�D_R"��k�$�両�Q\~��e<�Ϥ@|�A>�	)�,��5��g2�~*�I���D�瞫���j�V���������>9ՍR��߰��%��ʎ���02�C�����Mُ��ߡ��ˢ��΁��wq��I-�n�d�Wa�69��	D����-K�����E��q��Ap�<����f�S��W?C��~���~*�< ��	�6����� r���*8#����=N�t�*g��a�N���A���e=l�}�y��CW �m��yn�]���UM�OQ*&9�ǿ�q��Cv7�}W��,c�I"
����X�h��e��ot�ّ=�u[_5�`�B�����V:T��!��D��"w
��� �tr?����--�B�����1��{����d*�=�dԸ���HZrG�:�m�BJTI�nҾe��KȺ/:W���'�;Lv� L:��_�����n�����l�^&xe&=g�&-N� ���G	Lx6���T������ƵB}��-[���"�����+��\J��"�l jd�uS�_�X�cu��d���A��d�c����fA�Da2���'�r�5���8�\f��{yXY���= Z�~Xy[�5Se�Ĥ��o�P�.7���~�lHe�b�i���c|�ktg�>zzŸ����V҆k�O�'���^-s�ƽX9�#�l�*�[����Υ��

fl��
�Ė�?�/�����=�#6�wkY5'4�Ҷ��%��5���:�鞁r�& �q499?�:M:�q��"jJb"��1��EF�J�r���|��ŀ��'1�<-�w��؜2q�iO�4K������c���w[�ǘ�C�V@:���9_"��Ecc״����bK��������[���z_]�͗�l7���<�{�� �w�ǌ't`�i�r1�ѳa�l'׊qI�s�MI-d��12�,�u�=Ed��ђi�͸pq��b�����<F�����g%ŵ��O��?�A�u���~2I���V�h���G�c�k����N&��:�X6���s��@��A�bF�����cn����!�H���'�D�g��`}ExF�����nKI�"�FFݴ�3D���3�:}0�b�z�)Q�j�֍���ñkC���^i�
�ǰ�A��2Ϝ-��]�Q{�r�Sd��iG���n��OC��^7D6�Z��5ӄ�}͊w����ry�K�T������;�xVJ}�ll��8�O\�L�w���A{�+�H{fjP�;�+�$?w���>j%&%�*Ӓ���%�u������f�5a�շm��@�H�xll̻`9I�t����U����k��M�'�u�o��!�do��[)�W̽ON�\�15=��B�U�f�3�#u�L�
�z>nQO�B�=�>��M`h�-�5����ѿ\R�}1*����W��~zE��ӥ����E��-��y��m�v���:������;Z3���?>nD��]#��
ȩ���&����,xz$q�K�gO�E�h/��>R��l��:9��4u�191���{��������i|�9;����M�p�Zq��n`�J��+�q���*�e�l�ciJKKc���,#X=�Ӳ�!p�����'��Ƚ[�S�J���-�M�/�#X0�z��3M���L�5���$�Ϛ=ֆ�|z<o4��D��F>�LIV}�NTd��ǉ�B��L��6�H���]��M���㉿r0�;�]�"77��="��T:76�FyMLL����z���=���0n�B,EKG�O1֦cx�삠�����qvn.��2�%������g5�J�E�ʑ��i?&�=�o�6p�
�J`�������B6�.���c�����BB�Y�sXM��w�Qr�&���	��/M|C��MУJ�UeG��MN��]~'<���b���."0y��z���\�i_ff>BF_d��켶��fnn�>Q?�s�p{>���� G4��+Z�CR`L�v�4(���.�c��kkk��O�'����!M��kzu�91���bbb�q�#��*������ V䬦����N�!.��7D\@���2��I�N.�8�9U�	q�����t��e��\� �llƗ!���[���ϟUUDFՒ����7�r�1���{�����?T8�l�ZPw����Y8/:��n����ߡ�����&FF�ꞕ������ �= ,�&���%�A�˱�x㨘�8�|�E�$S�P�M}c��=����\�!��v&ϊ�����+'�^�\�¥�O��и1�+d�Ut�<���׸�Є�_м�2�^�(ڟ���-@�K~�5 �FH<����3����-��0���CLE��9}�\T��S�h�B����|BBB�bbD*&��(7��f������]7޴���Lk ��w���@���Ї�� K%��,����I4���Fsv�
;���N{ǯoo�u寨IܐX�~�}[fN�6WAP[s�D��Pi8z#�9'n_�o�~{��s���N��!�����RKG���@כ��e����>��K#6�4�ie�$����`_�'2y��/���^�y;{���͛7�a�;W�|�G���P��>/*n[��
��m/ �s�a+j�.�"�N��ǡ���Ӫ�[3S��cj�B����1F\�tsEVrH�]���1>ԍ�^Ou]]@�����[��åpOP4))�o����pT��i���~����`SSӨ6+��y���ݵ��|{s�r��( k'"	<�Dm�O@��БU�Mΐ���u} �ein~�'�T¦�J]�4��t�~��h�� �V��3�ǻx0X,�G����"��H�.�q�CF�y,��Àx[�?�c��>r233��Y������J$��0�X�]�(�Y�S2�0 t#0���V�%���E�4n�E�2����T���G�#5�Ͼ��?��'��TdT]���`���1�QD������
�Z�X��]M�2H���J�T�킮z~LD
��M����5��-e���^;d�mr�ɿ�.��JzU�B���ԼCJ���˿��p���]-P%�@+��]�9G���-C��%?)�(�"�nH�LY�g/~��wO��Y0�Ov{��{�/Ϲp��WC�ys:���:�mU��`���#G����7:PW�����?r����Ȋ�Ө��M�Ccݥ�[�5��| ��))(��u�Ƙ����-�eX��f�{��$ҩ'�2��1��J�srj�����zj�%�U��r��=��޺���YM��D_!�K��;�N�<<��Zn]}}��50���HaRS[Pԩ�q_��h�egow�ؒe�ae5"I��I������)��f�Aitv2L)g��ډ����}�o��"��u��1���$!�y�$�G��H���b�5S�]Y�M�íM�۷Gx{�nB[
�n�C�j���P�-��~�Cļ� 	���Mh#���[������ܹ��z	��Һ��M>��eVf2	[<@�Wij<522��5��R�y��{�@�цJ����z�F�E�8��@���?�,=�0��7�d�/MmN��cjA/;����2�hqG��S���J��>z��/����[ ze�� y(6�5��C8ڇ|0��s+T���S�k��������"c��ivP�@�g�.���N�s�n��;Mr+n�w���Nv`��z�'�٭w�r|�?����E�1_���Obr�7[1����#�۷o���& B�!
bu'�Y�<�DCMm�]� �6�st,��4��7���Ä�L�V��x\hZ@���˗S[�=.Wmpշ7N�tS���8����ٝT����6m�PV�M����ַ>�t�hɞ��j@�P�U?z��ᄀ���pj 4lq�{i$��CN8#d��X���Kʴ����Y;bKS���Cj�m��)����H�K&��>��[@+P�KO���H>Kk�@�s����!���o]��X����i�jԱZ�xxأ�.�B�CNK���DM���}�o��N�&�����13^��P4���d��}呚k��Aew�2���T�]�X���Dj	��+s�i�Fv�ͷ0�(����ଔz���������(�7+U=wK��(��?["��J��W�/Í��:B����w")�AF;�5�����J�,^��>�Vݠ�&��:��&'�ڮ��ȓh�T�K7e��k����Ԇ�<�ڣb]Yg����e��n#Mŗ��ًuwN>����^5�#+��.�8�x/GK5�uڢ�iӜ8'�v���m��2��ʴ�Mk)H�4���S9�&����w0 V@��,o�T������,|����$���:6��P3557����K=���yAs�[��qԽ(����kji�����zpȱ���J��.��~1h'��E���`wW&鸰z�ƓVVFb2ci����"����������kz&��s�[ȵ7�~��e�w����^ʳ�>/��� �� �B���&�TTa1N2�	���
66�������ή*i��Lbaaq���N�mjBX��~����Qp�YJ�}G��~�������xR����k���ׯ�y���"�yY�H';�L���2��L[988��z���/t�r�L#_�~���޲A���7�)�, �(�a��H��Xse췽�x �W�`�+��)�{{E���e�F}ikiYhyj�vȲ���7�t���j�&IpΔ]N �w�b�b\FZ�2)�_H�A��L��&�Z1��W	�-7>^P6x�FIz�G۫�/��VK|ЬGq$C��ec�z��v���
ɍ��Z rm�rRh�v�nm�M�h�˯�P�.�}(� PX���aڳNz����t�ŕ��2�
���?��2�Ҙ��^��2����j�;_t]c�Vbr�"�s��{��8:N�*��]E�[r�n!�9����"55n��ń��Yy�@陛��̚��g���,�����9�O�Bu.�C�Ά��I�$�I���z��6������n��D`HKD�.�� ����.�֩
���Ns�� ��V)�}{d
����tK�'[�k�x�+�4S[������*PN��w"�p�s�K1o�ۿ@����=�����Z�m6�����Y֝�7���E��L��ױuD���*h��>��અE� ��
4
����$�������h�g��Z�d$��u�'T���
l�Ҧ �ՑWs^n��cU�67��Ng�d!�L�5Ԑ(����<{="T̀D	wv�Ia�z�h⣃�1�p�*z��1G)�?al���8�F%�Ѵ��8���f�00�=�}�-""K=��+���k�xE>�G|���6�~��N�lh3�X�G�=mL�+B�l~��}��evv(�n�j�t����T,,,,���%�n���t�	1���7��X3g,�x94�Li�L� ہ���p��`6��L\F^�n�r�(	$�,p�jkh@M��ǘV6 ��\.L+;����4>��&�)�&�+Z���UUc�JO����6���l�� ��Dv�j�~��a`J׹�����?����~/�2��'j�M����Z��$5s��O��lc�4�!P�t�J���S���L@���h��a.�lZ��&��L�Z�88iXT�ӷ�E�S�p3��27�]����H�i(Jh���tV֝'����bL��:\:�L���w,�S���TTTȬ�"X)Q,{��0�
+�E�Z<���I��2�`J���o�t-�����P2?��i�U���"�0n�-)�![����� \��Ą]���M�6b�I�)4�n!U"��143;����XB��J�ejj��]`WK6�k_sች��WR��na2��#�#���0�5S��\�)��.S���a@ R9c��a�Q��`vww7L���\V��\���Yꠦ6���p�i?�ǎ7ͯ.���l�fں���J	�9�)|[Hi�����,�"��p ���e�(��?}���������2�00��I^��ؔ�W����WU��9!~օ�%Ւ���X"b �sT�����n�qw� �C
�k�ܜ�Dg�q0�d
���fT�Օi��u��)�*4���*p����� 3P\U��S$���6�J��a����S.�U���f��R� �.�����<g���^0��i���]��S�Z"��`)�B��d۠���D�*wF�#k����	� ih�2�7��MP�(=��F�a9�����TkI�7a^����f�Q��T �$��=��ʿ���m�����D���o ��q̏IèP��a�PM������=>�R��x���E���J�ؒX��\�2�M@�]pWq��2����Lʋ�O � HQ,��`i&=7�y˖-��f)�5.]r�K#�J�0v��r������W�hn�LII�#���55b&���->�����U#�0k~��+�Q$�uV���ٚX�+:��N��>gep#@y%$k�ǏgT�f�/@���9�@{́p�A�r��#j��j������x%%b[22������� ��%uu�Z�<�/d��c��DfZ�պ��-˿I/�j_:���JE��l���f*��t�����V��CϹ���=I�� �9ҌT���
h%���q�Tzf����3��5�o��7>��K�1�)82%(yN|���̀�ի��4J��]rJ�VCY�ꔔ�Ҭ�Ps���V�� �0zw>��=7�"��<e5�3u<Gr�a,������^~bDtG ;�?�829��R"�:��8fP�=Sc5������v@�]���K7��;����6�r��t����-\��0V�3@q�Z8<B��hqhhh��wS��m�N6<�[��Yz_�梁�_í�rҳU���%��ˬq�0�M~���Ĥ�S�=i��T0�N�ѻ�;������<�he� �����>1왮�eٜ��}�%*��o��%�aEg���x��T�P1��K����.dg��ڑ����.'��k�v�bM�o�Om1|�1��s���������R�3<����c�n�6d��I����Fl��JQPT,���|�3��s>���0�g�&o�4�h��秙p����d���X�����V0_Z�*����،��H�hA�D���΂���w��۾Yv9�˷�)2�8|�M8���.$�`g��Y�Lby����Υ&�����f�Xd��͎��ߟ���hLlF{�%T��a��1�_j��1u�c�ToqL���m�K��K6GY%Y?/��B�:-�;�y�^W��x��WeZeڢ�vxG�9�"�e0",��nT��5y��(��2LEؗ���QC��w%����1��O[,���Fs�M�S��j	���������F��[�����a��|����͛2-ڊ����؃^�$�.V��j��c��`A^̲C�㽕����������#��)������"@p���p�g��C{�2\O;}$�sN��d�d)#0���Z�?���RX��O'k=�ˇ�@RL���UKK�o]*�*�&��֥\*g�b��\�G؜����CK�T�C��:BRR,�}�'��u�j��'6��a��r�z��q�>ʂ����z��m���>���R�܋�|?�%QM�j�g�Z^�(+��㐿De�dZӗ/�����򳨑c2<����G#=.-�,��.�����@�e���VҲ43�?Y	C��"����mN��ab`�	��]��L���|I����Pؒ�����5]i&�Iꁵ9~��k���{|��^]C�Ǝ��J���>+�������)zyI�� -S�tN��L%n�����֝G�J��_љ�"��-����M�J�V�]֞��@�3�
f��I=9�?;��T��]d�1��(x�ºާ����U�N����R	Koa��3�L���Ց�����h�\����[i��ӳ��N���[̓���h�oh>���իW����M)��3���.d����R�"
�J��VV�ᄱ���|�������S��O>�:U�P�ѡ������#T_�����(��$��ob�� �Oc������p0(v�*�C>z ��S�-߄t-6�i�`f"Mp��&�,LU{E0B�#"��L���i�Z\S�g�3tr^QQ��"�!z]}pP����H��{��>�)0=kK씗�?�onn��͉�>�R߯�"��$,rW��)�.��R12�Yx[��o�fW�,�3�\R;L���4~�qgtt�ѣG��-�'|�2�������~___^A���ü��dӵА���E
���%��eZ��ӂ�ެ{������u���Ij;�C��s$F���5�7�,��$
n*bA�8W5��&'���rr�O�k�	j�DD�UOx��
&�UR@~Dx�T��JOW�����L�LYy�,���.��oE�����B�y����1	�a�J��/"�W�� c�{=���렄t�"ڎ�oǤ�i)~���0&�@�}������Rd�g3�Hi�Y����%��=?;{W��� UU����H����4������O�Y��e��{���U
�����VT"�&���&��h�����ՃW�ĸ�,�8���i@b+hWVY�?���:��Cg���������߿�cgy������5̣;gB�͹}�O�-4�i��7545�ה �ÏS5?;�Q����^7�5,���SO(*.>	Ѽm�L
�~c���f��B����k����>�lM'^P "ǥ�ӥk����D�s�	������8B@awτT�$;O"j�!nU�����*~E�4N�9� #6IUZY�j*jXu���Q4�f�b�ڈ�6�����Ϟ M#!!�Mz�4n�)b.#��LP2-�*�����5NI���rH8�2�wg��{ݐ���O�k"��s��J�N$�Tu��O���,p�9��GO�\�ؘ�职o�����s�;�kk^�sDn�dg7�v�O3O+�^\\��4rS+~�X��*.6���R.OWI��)�I���悮�/?ջU�?�,���֦TS�=C<o��뙹��W�?~�8U�*�N~#'�̮�IC]]�ʕ����g��]��J��5����Kt�F4O��@<�r����3�����1fM���>ȧV�,��SV;�ip;3�rB�>��%������Ԧ =(8X{�f��'��p�L�}��u���P:�f�QU���i3��S�)S	�7b�^F$���9iA�b�y�0�(����-�v��������m�?��������0�H���
��lS�MO7�ѣ4S�]� ��r��K��&A�x�t�޿iӦ #M`ZI�b�}����8<]��C��룁*�?-�!�Ѵ;��Ғ���/�¯߰ӥT��
�$ǝH��6f|R�}��eF��x@9$����L��c�v~�0 	�kKS9'���ܓ����{�!�8��һVݡPVQqP�6��! �U� ү����=�x�J���:6�8���
ŷw���aR�����ԚA���Ƕ$Eq��]��yKK���EEE�������������xq��	����MԲBBNk��v��D*R̈��W��ޙ����<�P^9�>���uu�ж�VR��+��	Dp�l r�[��)㌐h�_{�����\=�C���_����d%�C��!�:+G<��>�ߞj%�}{�s(;;;���ӓ����z�����ԡ&io+�'Y�������H������玄�C1#�� ��sr�ʍ�Q�#EћY8��ޗ��9T�ځk)�s�&D����8RU���U^VVXX(�9NP�O�1�755A�t��^���gv��wK�LrQ�Ӳ�����Х�6!{&�znn!l�����~H-?&��N�<����1I<�V~Ю=~��5J��s^k��F����j��vNR�����{�,'��e�ڇ���m_ߕ��@ٔ��ą_[%��|�u���ʍ ?���e��)�k��`e͕t��>] 1)��e``XW_�50x���$���<z�����±�k�C�}���f�oKBY�kX  .�ٶY<;�5�H��-!�^]=�`����x>��t�����/n&6��RV]]��ك?2F�o3�G�6�>#�VNNg�6^��&��#5p��&�~v� �>���?i�ʽw.��	�慄����:I��������@*�6�f흙�T�üm$��V��BR"{����6�&�B������4�b�萎�]$뱄sp8�뺟c�����y��<�s_���]��}������/Z�}�`$�8Ӌ�b�n8HZ���x��jV�ZB�B�$f����&Nv¡/2V��I&jn�p`P��l�V��c�(i��}�:tI�u�xAa�j�%ըY@�'V|~���a~X�d�ɿ�)��5���r��Iv�>��e˖(�m����c��}'0��n�A��yN��������ψ-��o�o�u�=��ْm�����8��>���5id�ΤC�{����K�'R�����h��X�V�3ˆƶ�S��~,a;*����{(�u�U���4�����Py8ef���nVz������==����?�8 _0���9i5��S���'&&>�3���nrWi��_���K�6��M�v9u[�nK���8�:;�0�g,�R��R��յ}��b�rM���;�-�לhѺ���z�ef���J6��Xl���fy�'�666G����#T��� ��&�������g���|6{�h�~M��;����R�w��B�4Z�@  >w�,��#	Uź�I�vj�5�y�z5<<��q����:S3�0��f���^P+�=�� �t'������AU���J�1�&��r,��*i��vv���iT��@�2��g�����vc&��w��3�T6���Ny2T>66Fw�R+�������EQ�-��ߎ�`WФ��!�K]]����Gj'�+{�˃؊����X۷oI��"��&VV��c�,��،����{f��Lm�]����R��S%�m�:456^����X�h]N��o5-*)n�25ՆB�D��v�\ڑ\o�O�D��ge�}���-��0'ҿ��N�B��M2�����;��} ���Wow ʄ.�e�am��k�8.Jm��l����u3�OQ8C�T�3=xv_���������ʌ<�@�/c��nx���(�]|r�����f�F��Ò�[6�0�̨��X�[h(z
>�V<+��p���3�l+%�y����g���ؑ��ST#v
���~۝1�ma-�A �9,({55�5i��.���5��?���a��
;��8ɚm߄?�(~����f��m]+����ג�&Fo��0ε/�{�uH��YyV��?��Ηa���7���Y��2��mtrr"
ǹ��iA�ܻ=~�s�Y+_��Q��㣘����['�p�@�]�wFY�&�9G� Q��ۉlH��n�dԍ(8��j�ؾ@Ȭ ��9U-]�^���h&)������S��ףYYX�OMM���8~7��l�~���Y��U�tOu�����L�x��!�k�[�M�B=9��l|�r�����_�R��Ԥm��7==�ʣ��Ԃ����;v�Αݾ}s���..۩���{��&�t��L��.ᄐ-�7d���Ǐ���\�&���[�BCCw�ݻw\|F��+���+��'F���>}��f�� dK���ZZ�����M�&���X��6�l�KJV��O�(�o���!�ܟ��S����-òb��{7�I������u>������|W�-��f��Op[y�����.,L��3�S����u�ЗPmQ�"<q��x�ν��[k�C{(R:v��t��ȹ�ؖJFE�������<pkE��������'����:��.BqyQo�'�X��x s�j>��u���ѝ�<����z���[C9����iCi����ᾀ�y��~~����ଐ*d������57�bM}��[�̋����'��NsF1���(*� )!)�5�U�P�Oo�el���@䫔�%Q�Gi�쁴E��B�>��ӊ����,���\��v������*))����Ԡg��!/���w�ާ[�^�r��ο?L��)P;!c�u��) %M�7Bо��]�_�|h>��S�y��<t��ϟ#-����[y��l���qډ�W��9V��bNYg��2̱0:�c��u��Q�s"���Xh
Lr�[��JF{�7E(�ǅ�.C��8;�6�A\] S;�� �v�]ٹV��7�v�3�^2V�h�� \�NZ u"6n;[[���:$kYq�(K
� W��*u���9� y�v�k�L��-j���y`���L�Ie���l�,VgM��F�=R�l�W�����i�Y���I���D��꾜�	�R��Tt��)3�� &8�f�'���h%( ?<�"���w$~hl<�v��9�U��?]<g{!��}H7���x�n7y������p��Ǐg@�T�{fA��.�^���)(q@��m�v)(�T��dL�u��1���Pzt���f�.*����=�K���] �&+����]k����޳g9���C��|{敶��	d�V�z�x�\e�=i��i�	�8�@7���Жܻ�&A|��Z?}
u�8�F����'��p>yAW�u7>>���$�[������~:8�����F��?����:X|@.��V�� ���>��j=,䊎} ��ay2릎�+��&�����Al�@�C�^i>~�x W�wU�r11������ؕ@~������P�ՇaD��0�p˅��ë��mV�UVB��o�lĉ�C�Tfϟ��8�mq������d�ȏy� ?<R�Y���F½{!�FG��������O5��SQq�*@p._0��88<�]nL��g�^��m<g蔯ع�}<��C�%�}�z�H�cU�O����v��HM�9O���q"�Dݱy̶���5��k��$({N��P�r�����\����ળ�����)+(W�#"#����4T"y͍N
M���(��W�]iS��k�o��������SM�1\�7�*���7O��O��a��Z��%�/���w�����.x�e��u�{��'졲 ����!��MUH2�J�ee{�{"B����wO�}BDB����䷝�=�q2��K@u�� -u��$)��3@< �s��?���)(��N*lĖ0��UhM�oR��'��IY����<���-C��޾�3���]"�����jh0"1��S�$�������+��u�[�����A��H�%I� ��/���Ќ�d��e)���/��+�Ml����#��(���B̢��5\�Z;s1nu �����������_kcc#4��(�2J(��
lQB��sM��B������Wp��I�]�A3�����is��'�k��C��4�|R�.��)���/_>���d��)�</��|A^�2�����*�+Q�vΥ-�\w~�'�[=p�g�sg�p�1ߞ�XұDMN�X1������ˤ|��P�����w�o�?���͒�[�
���j��]�D������B�=��7��[殺���P���?��o�K�|'!A&M�0�����>�9 ���s�)5�칧����W
�4h��A�zgGGi###���Y^�V���'Z~�A�R�w�=�ԥбu�� '�)ħ��Un���a~�֭d_��|S��^�9���C���Xjoo�fL}�_-!���.��O�*��]b��f`` �}0���+CjU���ҿ�f��nhI�{�r���K=��8YvN.���u��b����P����k�Q�TpU?��[�{���e�r����\�<�;��qTpg�	5xx��/�d	�����w �&&&px���y�C��$1`l�&\�ȉϮ�����nSH?RkKK��opŻ�]x�jk-�v����'�-�U��"�Jq����ɵ��~��]�eoȼ�-<9�c����P$pK�����PڡE��4gh�~c[ܵb��h��K�n>��������Ez�ڵ��g����[Ma)WU�4� �K]�Xߌ���C:Z�Aq���s	�o0�@���06���?}ؤT3L��o���+ZZne��v�
���FO7��Y��~��N%ԃ���y�j����q.�{�66t�>�^���mm;H��P�i���w� �]\W2��c�D�?���Ķ��E��C�ԃ�_�p-��ݽ��ҡʣ�Rf ʾB`xx��3e��frҷ"���gggg���y�����x&�խ������A���7}��Y���T�Ì95P�F��UQ�1ϗ��G��X�jUگ���������6����8��#��AT�?]S.+(+[\DJ���s�<�f��9x�ch2��O�/�gA��_f��qؤ�o]Od�AQ8�.̀"�*�i�I���*��
���LIU�SΝ`[�*@�Wc����ar&K�@P�1�>|8�����6��3�Fr
�ъ��}I���N�;�������㎊�5�s��Z~@e۳���K>�ؕ �Ѯ*�1?(O�)�b�B���r�Q�[{yɃa�����\-j-{}�F89wi�24���\.��;a{��`:�(�G�5Y���u��d�DF3ù�Om���ۄ�5�ɉ���:���@>��wt�'W�}�
�]`�˗/wd����]h[;�{aeݔ��\�g ]	�7����OL�(�/1�b�����4n��0UW�~b�����m�i��jrR	F�r��b���H|��a��ڙ`_ʇ��@��� D�YKHJ�*��5��슄Qw��[��d)�n���_/U��&�Ru%�K.�@���p&�5p���*�w9�@xd(�h�4�)��� $�#�}�W�.Ⱥ������mi��-IձM�m��Ȼ�$]]w e��X�PA̐"E�%#����v:'dfr�.��Ɩ� ��J�ob�� �Ҹ�q����(���LN�mk����_@���N�x�	�v�O��������>�J\Y򡇂9-���{�؀�Y>����#�����JY���t�8��Ą��}�p��m`bZOI�0Q��������=$���Y����۴�j{�^�.W�*\��AU�����4��ax����1|r�Ņ;�������MV�ώ� ������<;��d��� �E'����ӧ��=9�����.y[笠��
���Nô�{W�o��t2�	6����ND�S:ݒ� ��:���t�һ~����瞞�&3ї������^d@K(���F0� �<�m�j(���<�L�[���n�5#�1"�mK��u��^�����;r̝�֎Bp_@����秱 ����%""�K��3_�-�ժ� �}L�Н��[�:���3��UubG���~ZXx�t����
Z��nL�Jd#��!|q�To�z�8<鉌�f���R���>�(kTn\��m�1~n�;����e���wC�K
��
���\	�`v2\;mt���ӚA�V�O���������DuL����.U�{O��!��%$b���"���ܳ�ϟ?qL���p�V>?�@�_m(�̱ml#c�O�6�Ӏ����!�i(��;����Y,Ǚ�"!W1O9������3�ROs *��66���x�>d�,YEE�,|R���X���,q?DzI%����'>�Uu�$��s�������쟮j��d���P�!�Gvיִ�	,h� �@%AmR��6w`K%q*g�����k����4�3d����EOk� 2d� ��Y~Z��,�Ť.���bZ#!	��ӈy�l�J����4V�'�1��O��z�}��o$�J��#�����h1�,c+��)X�3����R�&a :Ys�/�pe�Ț�?��0��y{��-�����砦�Z�$A���4�c�ɡ3�xC#�]0�!_������ �4�2�i�e��N���U���9���j!� ��F!����!��>����Q2��|3L]���'@jڒ�� Oo�V>:35��_b��EAi�D���)�P���x+�W�Z�z<�v+=�چ�=�nBC����3�J"ԧ���3_�+;�H��wvn�w�m4�L�
f��� ��?���ѡ����ں=[���)l����^�v�H��4��,����95hB�9j{��" �TXI+[@�W��~�6�@��`�i�喰��ɦ"�	�wA�l�$R���ԟM�IU�*e��vZERJ�}g�z���w�b����9�o��ï�#���$p �d �
{��!M,��8Z�.p��=�����8(Z�E�~��{D戄L<kS���{�c��r���pi�]?�ɬ*nV����~$�}! S���TO��fPh˼ǝ�	��f�]O���i.}Z��0aU�Bs����k{��hU����;! L�<ht~UWg@]HEx!��8�b��FB�qR���i"�ʄ^]λ���CXBңlM��*&�!	s}	���Ɍ5b�_���	��xԊA�B�Ī���h'���*���;�,,�O��Y��f'�r�3N�g�^��O��/����ȭt� ��z��V��m��BWo������7��s�]�"�Un��_4���ׯk������̔���$����߆#���hM�Ђl�S�{��a)�Pѻ�~W����7{3k�hO�4��M~��A7��jTand�E��" �	:�l������p�G�h�㸋|�ր�߭���뙙��r���pÛ�ܓ����u�m���B0�dښ��t�0�\�����d��q��ʵ���x�S	�%}�\����e8��Fk�=UC>�,���U_�O#o��������b�ƍH]M䘷��	�fL���n:r��
q|�8_��P���*��Ʉ�$>�Y���Vr�[;r����(ܰm(-���¯<L��ʎ���E�]#Nd�y���6&��e��ŀ�?AM�f�/_��Q�)�]]���$N��A|�E""�޳���OG��ʷ�OzJ��fn�rhȵ9l0�X�f7t�1{{ϱi�}�]Ǩ+eePN9^�wj �d`q�b=y2�q5���3��a2Q,��ب�q,\���c!�o)�s���օm3ιw��v����,�����v8I�!���#��]���/��Z�<(�p�������)Q"2QxzH��8a$P�5W�E�&(����Js��k�&�ʹ��^��	��޽K�K�@:Q�@�eEǜqsۉ�=Zۧ�O�8�>�f��B�
!W�;��~���������t���L�K!j��kntm-;�xţ��K�^������!��ρ���eU��lz��B�nI߹�#F�.�#���ߗZF���E>�m�N� ro����ݛ�(:Na�fg2�w��f��;2��yʨ�9Z%"99����%M-��8���J����8��oX�pa�caS�=e�C�v �Z1�pP�T�&H��π���ϨMi��W���s@��c+�R"@�@�r	PPRZ�Z	{�8�/�]tf&����EWg���l'�ߤ�X�r6���NkL��O��oo�%���� ķ��s��S���^��i�v����|�����8�5�=���T'�����Uu�)::����l�X�
��]��e����嗀y���AZ��h��a���<��`Hdeq��=ggO(Օ�p�͙3�*[	*�jjk�!q�%[�V���Lyɇ|�Ɏw&7۬[����)@AEe�|tFom���{V�Z������>�����MćJNǝ�Q8�r���}�$j��n�z9�����m�Ǭ��+3+v}��_�3׸�U��j�s,j�"�"�C���0!��v������*+�X�`)ǋP� �4��7t6��Ђr��e�T��o���X�	�4a��=	p}�Z�57�:�R��H��8|�$T��SSSw)*;^� �����j�g��8"�M~�SRR:��k�R�$5<��#��5s�w|�����ޥ)�3�\	�g7�b����d�>/*@Sg�#Sm��S�i��8]8�70��Z�N쎗�=	�����8��x8F��"U+�,n����� Q��[	4���G�p�ٍ������M{���#u2�)ː�r�#v�����!ǎ��<���B�s����4�X�JY�%9��
v�l3۪�E�_ ���Z��	�uT���kϱ(_	�pO��,�c�.�*��4ྜ��$����P�,�� �Q��p�̅[ 9�`�����+� �]{��x#��	.����U:�F\<Y \��X��=��$����`���;⻁)"OT:����S��H!qj-���|Z����^�V�����遗��Rě��Y��o����9�g��\���EQ��k��$%�*kB��j�,�fL0�d,�a쁘�knl���lNtqv~�](BVR:E�8�yy~���{ÿ�����FqߟA)[�ؙx�F6�ő'KYJ������[�4�ݻ4���ň!��Q��P�׀Q_�h(u���k��9����n�sju%���������߹s5C?��T���w9;�b�2vO�币\5�"����'�{�4�q�_T���j��Ʌ����<xW���@�27�!ܰ�2���fj�՗/_�z�~=6G��wt����!����1��7{��#
T�i���c
e��t����"��HE+�MT]��BZYӼ�{{�].���Bu���N���$Q|��Wu��*�NUf�"�x��U�ȍ��{Q�7f�+�������5'�1�ٞt��"���A�)z��>�!ssz`� .u��%XOP�Y���z���rV�������߉F�}'��}[��Wc����#Qy���7��s۰xѢ����[yEv^{���E���I+�znn?��wab����WZf�:�*qK�G\�F��5�}��wAC;��-Z��3<����R��kr�6X5&��\K�l��G��GFܨr�@E�.=#���.}p�.55q$Q��@�y*H_��ĕ��]��d��nMMMA����g�����"l;;�N�5�i%9Drv�,�zP����Pb�A��2�1�J�(GjF����.�S���	�6�p���u�7��N���T���4�j�b���FQ��o/^īh�͘�"��[E�@��m�k�Y��~����X�h��W
��8������Qltܒ�3��>���-Q���t��h�F�ZPY֔�n��	[�b�D����ڎ���Hq�~�.
DP���֐�ҥp�ƞ='�o���!<�o�eq���̕H���q����{��B:N���c�&��mj�	�Ŵ��I��]��}��]�Ꚑv%3Qh�9j�D��t�O\8�%IEsS%28}���k)�p�~M�T2�r�G�Jx���,�یՉ*ӑ}oWj�Ml�!rr���zAb����x�x�;4�C�A8�9RQ�7Q�Bn2o�L}���9c���ca��O49����mC]2ؘ�M���m'��t�C:���G!�\N3T�իSSS%>Ö��&1�	j�I��\��gPt���*��F $�GU�=��Vq:_��Ã��:��m��x��t�Gƪy����_����q�im7��Ӻ�J�o�k��|{f���d���ݻ}�
H�4��(�#�}|�� hi��0/�U%i@���������])� �����f����>�]$&��*���j�7
���AK�B�K}=����gFP.�"�;��f�T����f��WVV٣�E�7��k�.���6Ȝ�é��K�8E_���s��J�䁒�s/"�N~�K]?hݦcK����p��9?�%?�߿62B�D��?}�
���y��P�AD�⡇�-��n'�ɓQ.h	�]��
�m�J���6im�o�ݚW��^���㟗ѳ_�0#������A��s�o���̞��>�5t�w�ܑ�@�12u'.�ӡ����p"�d����DBY>l_:���-̷�#n�y�;Ed��l�sJ���|�v^* p�RP��(S��9�c�ri�#�4����5��x^�£JԒ`O��VT�t����l�F��V�G@è����j�i	��������$YP :O���]��bRL���7lW�e�Z#fstH��*n�CzJ��u�&��3��7�𗊦"Ui���)H ��|{ �zV`�8�*��4��xw�
��gLŋK:��߼�����-X�ҿ4Q�..6�&��г�����vws��:��mIT�[v$j:KԦk�>C/��3�#�T����QAȡ0���X����'�_UU)���f5��3�%�3{����H��"�fRd���f�;	�����������}@�귔ym�{߸zu�ڵ�!zZ�����/�s�՝Ri8��uɒ%��xqhf���-�6�VM]V�z��MGp��f������Ȕ����|*�����g����+：�	�P2L�3+ܙ����dfŪ�/�T�`���\鬔��?!PxfZԦ��?"����K
��qp��q"5�!,�L5U�����66:(�ɉ�Z1"���9�EDp�a���~+"c/oy��hNy�1�6���;i�ˁHhN�����O�d�,ߔ[0��<��� �ɿ�>����A����l�BQ��������Dko�����CBu<&;إ�aɓk�v@[٥�n�}���)����c�%]�J#��Z�ۚ8�hZ�����O
�è�~;;L��`���B�C�pjQ�;jMq#>))r����2!LM���.�<��]8N[���5�F
E��!e���*|�.UU|*z�2}��<�{��J�'{Ī9����79��B�Ju�k��chGmB�l��Z����(����]k�l CaE��)>.�?+Û�-!�o�Z!ur�5y�3CЫ�5��H������
E$�n����g�k��Ar7	R�U���h7�'�R33������h":����rMJ�=���9ei��R���p(�z5H�U	z�Mėr [�KC�F��n��(�}��ɓ�.��u���Y�TB�!��	���~`F�
:�f��i�WD���|> �օy^��K�.�X�i(Y.��$WQ�5��F oh���*2�tHi3O��65��/��%����{�?~�Hɉk�:�>�q�m�H���1U���z�\�u���� v�&�M�FI��X��u� g���5h���5��q�9~���Sb}�����B}CH��[�d��/�q��&U+�@�p��gIj�)\���:��)V��*�ѱER�"N�E�5~���d�_���{�Se�����K]����=�uߑ��'�v�-9�ä�N�c�Z�۷�����-�� ��}�sM��H�󑓱�a�D	IL��Lq;���PBth�+�S��s'>>�U;n�u��t��3�����h{��MЎ_:���Dʽ9�V�-X'V˨a-���+��k4h���c�Q��	�.�<��s��q"6�D��S��."Nq�%El�MG��c���K�����Bh��Y�q�UҥF�8x�ࢨ�`��]��6	��<߈駨ج�A$�Pх� �w>�3'�?�%]�BBǸ�݋�����/G�����(����v3�5@]���D��G��G2a4�56����
��񧥥|��q���з�
-k�c�MNN�/ŀ�Ƈ�@~h�n'�����.�X�Z���]2,��z�Ğ����\��#Q(�dddn�>�&8#u^�ג���?�J�����1�T]_���w��s�O���� �7oR6�b�����^'�:��N�Z��#�P���LЭ�ˬ���.�.M�n�o�d����b��EkW��n�����a7oB�����.,#Mu�08���8Fpd�C,k~όq"���5@�T�Q���Ή���knlhh�>}�����$�(h溺��ˣ��6\�2��4u�l���6��h�o��%wsA��&�N�f�s	��PK���V'2�̈ ����.�G�)v+ձ�\%�r�&p�8����Sff'�����ֻ��5���3����p�����C��J�{�q���֖�sr�!��	�T"K��(qN!Hve�i���0V�����ܾ����G'�����)a�o�Z����G������&�T⿨�����~�������U`	��U.�8j=a׮�x-c^L��Ν?��ݻ��혣�xn����b5v�����X������wD����'ף-H+�o�Ɨ!�3(x$�Y�.����6���f�����R���R�;����CC����Ū�S牐��{�������sr^e�Ƞ�|f5փ�j��������fq�[��R��ǖ�gMґ�ܾ��?4�StŷX�Cm\�g�|������	�|���Th���}vz""_��&9����aj�)R���b<��>C?�x_n�j�s�b�24 l�0 �T�L�Ω�w�T@�'�G^�+O���-���^����kD��{#�����>�G�@�-�t��X88����~��5B�q��_�6���kB���>|� ���@VW��I�^ F)�j��HJh$�y�U�JR\:��a����B����5N_l���J5R3Հ
�O������?�����2Nx?r�������(ť��t߀�N,}'��p�xg��VXJ��=���Q��~�dv���lE�QE�TG\�]�@�&E<�E�֯_o�J�[;Z-�xj�9�RZ�7ć������G�l1�z�nS��7�j,^��H��a�z=|�.�tH�:��D\��e�޺uKU�e����M���#Y�����+�.�gB͘�iv�Ӝ[�&gM�3`<��[[[I	y�K��k,��3�_���'�j�u���Z[-?��:�M��|݋���+4u��j?"d��S��	m�.Lp#�u	�˸��}jj*τ%��]T���˺u��恎C��k�*��^N���S��N�ݱ�\�i6WxѲ�GDQHR�	n�|�D@;�`:��|�c!X��V8wy��O~� �]�o�ћ�i��U�����[C!�͔P�n�kǋW�4!B�bi�x��̤���=����nʭ���6+>A���&1/��9��EB0��;pI�{�r��}A�P�e$�Ɂs�f8}%<����O���i��+�/Bb-d�v��W91��9�����!P��
�F�k��l<������"!	]-.>�ok������'?��j/#I�>xff�xF�[�.�DC:��S���t(.��Ҳ���+Ҭ+��{�#��0q�bݿ�wW�LU2�u�ĉс\��y«���E� .�t�F�X�&�fdfZ��L~�]��KA�Ҙ ��klFi��0���&��b�`�ڜ;����>0��f���!||�CO�:��@�[V������o�i�43df$�<�E%2;;'���㩄Tp��W̦#3�<���qF]H�6Z�{V�1���!s�s ��#Q���R�_�L��e�\����(� �(20�8)(+qr�p2�����QF��ܻ^�/��2�4�vp�J�4T�� ��}y�X8I��0
��������E��Һ:::.!�V5m���'����Em��j�ά���B"�ԺS�j@QUf�	�s[e Y!$d�Pږ|�߆:�
�3�<�1�5��BVy��u囲k��� �#fꚔ�p�*d��V�D�к���cۻ$�9��M��sP����q��#��[ը�L��1(���m�S�J��&)�Vk��L:���Z�=�x��27��i���		ھ������H��\��ƾr�J�95 r������J3�>45]7�bq�xYV������ގ�ڕ*Y^`�|"C�%v�ŋ��aЌ/?�I��,���(�K�koV7�t�fq����K�'z1N^��_�K�T�)�?�(��}N0�ZLl��d|�#T"��ŋ#��4cl���D%&�swB.q�F텲p�
0����(OP���״��m�g��c�������j�T�[��w�_��N�$�
xZ^��u���V�Nb���!]}}���QA�,��9-h�F�%�`�Bf�$��  q�S��7{��<����e.�לhUz~s�Tw,�RU��JHU��}6��l&�_ ��ԩSWKKK�R�;�;'<3Z�����Sl�� ��vT �D4x�6?&��2޵sgm��V(��==�O���C�|��C#��g�eC����ތGH����9A��Uf� �c!p�-n,Y��W��2��V�������
 q�~3�z߽;�F�~	�L����q�rn�j�鬉�wB�kK�R���2������(�l��_T�*?��C.ke�5���$��ZZ ���p����1u������^uj�R��Z{��tv��L�)����M��<�'S�|�#4��7C0�dی����8Q�W�v,8�����ƍ�b��p�zzb�r)�io�Pl��
݊�c�C���I������>�R)h��!�� �����T���c4���DՁG/�}iE�S��Ӎ�\�_AV�f�L���qsۉ��l�����$̰�0�%��I��k�UEZ�!�+�2hm%@�}�;�[��oܹ Ҥw��cv�={6oh{���Z"2�^r���@	:::d)/5������C�A����
������
�(C�mp�yfz w׾}M�Uh]9���~�	d�q
c�~�^�M8cS�7fg�WA���&�(�����z'�B���ljr�s��ZZ�	D�ײ!����7���<<�d�`<�-�.�~#�t�#���p8��sA�`��k��<b�?�1Հ>���!	]EX����"U��a&�V-�T�pǕ�_inq5����ߓ����Ɋ�n�T�F�ڵ��n�Ƥ�\�q���n�,hQSU�cz��-m`"ll�*��}
�3�v@A�^��v/��>�d�d��G�E�{�����LN�%�����(��~qI�b�C"�N@(�/�d�������jM��)�z�.��ڬγ��%˾�jxy�F����C�7��ǥ�����V$>j��$O�Xy�rlOg�����Ws�s��J��{b�9������5Į�F��v�D��Dل�KL� h`|�3e�ЭsVH<'����Av�"	�j����;^��Ƶ�a�	|�	G~~��=�0ҟ?Y�,�.7����Xd;��MCN�K²�2�/��n�A����3�s_��J��J8��Ͼ�3��gB��u6�S�RL���ԙcW'ck��m���Y�d�k���� ���B��Y�f�R��99� 8�U˄6�n�$sy����X��7q���FZ�-��A�Q`�"܋�Rt��n�x������@��M��D�P�b���%K����� H�5A��ɪ��Y�|)ܞ♅yG-ɵ�l�'� �_���3*��3q�i~��nE�Z����%�xd	�[� O��-�Į�����U畗�u�����Z�Bk��r@w�7n��n�읗쑨;��5:�������f��6] �7˘�N������Υ �L%�M]B�v|�������BSUn�p&�ckk8�O�D�q�:��퉻�*ב��2�M����:>���
7���"����7�"�?CB
�mM�]\PL&%EA'\= ����FҡJ-���h�׌�:kW��mW�nI�X憸q9+�2�j�qI���,��d�gB�0QWiE��_��� �6�A�ٽ�hv.�2��j</oT��9�2���Ep�o�1�匰�	���О,���TE�#�LB)GN��������M$�BO셸�P�6�x�1mI�Ԟ8����)�ە��j�����)3��S�Rd�Q��p�3��Q��W8��iǯ�-����&U��8ea��-(��ړ�Í��׬�2Sr���5�+��y�H�L�܈N/]#��f���?�Rջ��L�)(���ڀ�q%�(�c����<ɤv#���t��|(��A)�R�$��T�F���ف�5�6�~c8�"�� �$��u�4��u
��'\�����N�7$�y�������E�)W&�py
�Q#�V"�U�4N䎿!I�Y�����E���d� |����xr^H4��w�5�Z2!����u��i8��<��ׅ�o��F�����'��\=r��%!�Q x��M�pG9�7�W��Ȱ̭�H�b�~���^P�-/�b�ƍ��s��x��wB�#ʶ
	���@�:�N���ϡ���ȴ�������m�ۄ�,k�X�?��F���N��<wF:aNkn"&5ۧ�m�Kh�Ϟ}����ˊ�Q��z[���h4Y�!1�Z�B�ş������o���,E��E)e���.Њp<�z�9�O�	��60�"鮉=p'�)�`@M��Z$��1�@�wB�q����߄=p���9I�<jg��X��z _[��s�O���x�h�dh����ʃ��!YYA-�r����9�+��X������
ߧU�4� 111��{A(1B���c�0B�3=�Us����A%�Rhx�b�L��.A_���R>����Xx8�SjN<q�`8�W�}��Bכ1<+�?���>�hH��՞�{�O��7m�������&&�W��(�oO�g�����f��c�<�U����fѫW��s�*F��<����1m���N���������C�U?~gQ�k�ѭ�孠�C�m�"�����*Jp�a��[��7�ڰ�g(J����M�%��V�kN�G~�����S�L�y'��lM�h���I�t������.b�}i���h�F��T���絽����G�|�hAǽ��/A_�8��ʖ-[D�^��2e}��Ny�ʰ���!��???f~�����t��~��2r ��1����Fg#�,�Xgu�V3WZ�pm�$\�w5e����i�A�F������o�4��f��	xe��)��A�L��(t�2O������{�1�%���eH)b�e��\����N�ŋ_�^p�kw=��K_��pN���Cp�eXX؁ȱ���z�V�L�̚ǜ�����H���57%�>;�����3zV���E����GF�����.���3�6�ˁ�����H�_�Z_X��(R+˘I��i|Q���a81��B����r�w����}<g�Q��e��{��}9��љ|�0H��U]"ɇ-��1��uk���)��d_�;��׽�C�>���⪏��37�jErU�I��]����67p?~<3�-f���ha�|%h-��gJ���V�J�,P���+
l+M_}����-�m:*�l��#�XAk��l�<T�zµyLdWz�r���
x$몒V��A�6�[�����gV������q'��-P���	�K�� �ٓJ��Y0�+m��L+�~M�������KbO|i����2vqi����'n;+]�ƳVY&������{��r��Kǥ�������[R1?e�G�}�����ܜE��?���d˂�P\j3�P3<�'/�4g[;/��Sz��x�!��'�`���3��C,�y|u��WNY�����ȭc����������6+�hȾ_�'?��?�P��3����2���ZN�W��
�D�@���}������V_I��3 �C��> �`aԙ�k׭;!����:���K�}�&��{������T���4E�E�	��*�[��ݺ'��m[ن;b}*%Z!۲��_���lZV7�U�⿵{���ѹ��K
���1/�#_qt�=��i�������S�K|�z$S�}{�O7g��6T��gܪ4��,-������_��}����eDF��v�G)B/Q%���֢�ۅ�!ML#� h�;VZ��ip텠 	f���5�c*wӏƍ,E�|�vZ�t��6������n��ILZ_�CZ}�}���e���E)�8 	�������^Tu�m��V���~VV@ℊ~��F���m|��@Gq���X� bҵ�d�����o���ɋE�i�\��d����^��)��߀j���2⒒�` j�*VU�{��x��e=�G7�z�sQc���;զ�A�e_T�S�$J@�>��ߴi�s�7L�)�Y!���_����z�x�JNWWO��ae�c�(����Q͹Q��d���a�1h����|hy2:x'�-�K'g��%�uRz�s�>��+�����c���)�6�šϑU���KB����CT�]�ee��â�AU��Bշ�tO �AL��y�ZU���
�8�v#*�X"5�/�	��lVCC�9�ut������'>�{��9`�cR��ѽ�oa���B����V���ϣj������ ��Bc�Q�H���,�9�Ue>�%�Ӝ=��q5� �t�X�0�C8��7�����Omz�ۜ�2��5�d7/�a��/���XYl�#P%2c����b����P:O&�!��b�Sqf��T	r|�Q}CCC�ݥ���-I/ܰt20Y����m��(���H1곹�������GfŮ}\N�XqMk��xBR%eee=S���6{��g�c֩[�	��lᘊ����#�������cd�����%�5{����5�͚��Y�l��
��Ȫ	�
x.S�Ͷ掎���9WW=$�9���B�h��<��!���!N������H�U��-������h���ր�D(eF��?�\2?�%��Ӟ�����j-�AZD]�r�4�>'����b�'�d�f�ɓ���X��_�8)��XWTT�ɯm�������z�}j�М���:���¥߄����t��珏��c�x,�/�1�9V|�m5 �)O��*4սr�"�5W�
�
9�������WN��wԷ«/��58������[ /х���׿���*9E�pߩ�]��c�����O��ޘ���~B����De~����S ����9������YOy�L##O�HJ���H��g��Y�,qnn k`Ph���..$�I��XƌF��U�0�<�G�8A�E&�z.�c��1����p��c�9{tO�ٳ���N�}�
r�{�����r�fP����~i�ˢ������~|�67�"Lc��7o�$���]�]o!�6"xϝ�0nsP`{A����P���W�1A���GG�~`gg7��0�Я"ө�����5;'��M���+{9;�#��VO�ܧѧ4��?p�n~��%ɸ�  �]݉;���l�>��\�U;̏)Ļ�s�⺔�jk��g�s�|VE@�����غT-� ��wo����c|����+�q:m��� ����Qq�!��X|͛U��R�8���rx.��5�J��~}do��y�"�c#h�{{=4���P� k7��\��4�����g���$�X�ӷ����q)"�m��C�Q�v��#9t�{ 8$$��IA���ƛ]�ܔC5Qy��JX���o�ud��h*t2��X� ��鯥ش��'	�%�ss��xA 5�����-���ܛ9z�;������c".~~��EdF$u'�_�#w�Ki�{�o@���'����kM�~���t���é)� >����V�f�1	�/��I��ҩ��g^�U�y?6�O���u�I�)�O?��
�?ܽ�f�E�Ϋ���
K���C��G���L--!I"�,z~��)T�L���:�;^{�Z03��6T����[��d�}�����p���i)�3�f���䕕��3�%���@7�u�V�"U*
��/�?:��i�ZJ�������0��t�2;`��i*TMb{u��/�ʔ�5�?�U���Te9@�UE��ҁ^^^�jN1�
T�mmm�H�P�-���0���{Z˼t~��'�r��c`�N�81=T>\PQQ�3�Y�֭wP�Ba{����a�,d�caS�~��7�T��g�]}�\ܾ�_�a��`c� 
����e�Sy


��C�8+�1ؕ��9A�\=4�f��n�Y��bv匜W��%c1���H3X�Rs��㍣�`��j��}��V����;���w��2����V���V:lN�%Q��RQ���19��Oٲ�!$!4&�!��(E���`0���<����P����������_�l�������������� ��tu	��M�j9=9=33���F��?է(2*9�C�F� �A	C���[5.��Θ��vd��?_f�}���f
����*�U^ً|w��}�w��'e���*��4����weҎVz�8xTI�y�zd�9Pe�AUƹOh�R^z�I?�3�-���4�� _�ŗb�?��xb�
q*jƠ�41���UWGq�ψ՚z�'00�TJ!̆��1c�Ur�A�J$7k�7�«�C��xj��U�'��Q�6��-�toA(�����Ը^%��I)�Y_OO2Հw5g2�Vr�'�*�ׯ�C����j���m�74ըI��.�3�T�Ȍt�X�I4�[n�H��_}h���h���
vZΝ2�������+���m>~~t�&�úk���uq{9`�Y{��C�������A<�mm�=а $�F���Ǐi.��!Q���������<
��.�<!���aRS�������L��R`�a�8nա�lY!��(�m����-Q���Q�U��BX
�Z��%�@���RZE��R�՛Y�_��Ga2�ȥ��rroBNp��w��,(���y�	�B��Z�D��>�?��I
�(���u[*H��}�US��]�������*�GJ,��N�<8�Z�z��2�����fK��|3����Ej�FY҇�G�G	��	d`���R�b��y�!�[�1�x�NUj�Z��y�'���9q�2�UP ��H�*4x|��άf���8@|�Ai�Q�l�i]�؂�f)��ԃf]I�xz>�;y}��Ǒ-kx�����6N��Of2��f�kv��d�k�A��r Q��Z�������B��zȂ�Ѓ�7�6���
�"�Zi.�e������Ku��K�.�c�X�h[K`���ONNV�d� � G�f�Չ^�<���`���p��� ��䙠��s�/���e���H� R�h����%$�0�N�����b@a�W� 8t��v��s��(�����@U�L�����8 �U��C_ݙzR-�x!�2J+Xʳ�!�'ԽE�|#,�)��Z ����~!>)!�2iot-ѧ"�e'۬)m����0Z0['2� ��]���j7k�KQ���j���ՏQ��,��;'TBJ�E5\H�`K:nd�_J�U	��}�Ŷ$PL����(�(j��%4�'�v ���(��s�k���P��?&A :C%���>}Zߖ\j����\y�2�Zmmm3�Y�FY�N�C2�TaSס�C� n>%�5����*p]of��������n�V�:��ф�ڪ�Z�¡� �<xpx�>��/�P�-����wC't�h�Bm��J,�R+q�$�
��Lp�({��-a��enn��&2����G��گD�_���ylU����t ��@��sh�������<�������bb�5Q��J��}uq����s��N�}����3�"Б�ѧ�:Zeh¥��6!�}�H韯e ��P ��<��R~˪��i_�F<�ؤ�~��i������2jc��TZ�-�������P��~��L����a��O�8 5�S�F�ŝvS%UU�`֠ܬ: f��N�R���d�]�B�����N̨�h��׍��6�Y5��x'Zw�X� {����e��o�n ��}��]�!X�s1쭲��/c�/�+(E�:��o���u:�6��t���4��&��3
E�x�)$���D强��k?[YE� ���@kL͍�&���4ܵ�݅����D,�WPȆ.A�B��c����F��F:�Ç���H�,��L@4�9�zS���C>�Gj����[���.��{���7o�xg��m:	J����jU��X��P:��{�O����s�?�EB�@���k��}fFZ���*
����A� ~b?Y�ȇr�M���Z�AYu����Yn۶Q� �,4̤6��9C����W�`��U-����{�S��+���r<�D�rz~0a1P�CY3f�م�H뻄k����9����)�����˒|�6�d6=7�=�vXkσ��gV��sj"���^�j�{~;+��5h�V(����D�lNe���J<��1C�%��ܩ�����2��RQ�]�Zv��ս��SuŌ��v[+ެ��L�ooGLS])�l�̞m�s�nDD��'y/<��f�/L�^�����?3ܐ��|��ͤ�w����D.)�w�����X5��nr`��ީ��p�n���ǪJ�KÑ��Y�DL�`���_-9��795���۷7cpW����6�?VI�g��H:**j?��V�%��Ol�y]����h�����"u###�ih�|d���2�����	�1cjH��U�^�sYs]9
�T�C�{��ڵS '���~�V� pn�c8D��k��J��ܳ�"� �nܸ87~P���:0��6��Y���2T64P�l�����`՘���m"�ܞ��&�ƧK�!Ս����/�srJ�	@�;����U����5P:1"���tM��g!�Ŧaˌ���/���el�/ P\��zzH�iq�����1T�ݭ���GF>�XE�������j���PN���V�0���y�NE�2޽�|���if^~�������Ix6#��`������.�a�7����tF�x¿��q���:�%>��t�1@�D#]S�R��b�jhp=��Y�q�RՇ@� ����8��<T8�|@`4X��k\^yy����3�P'����g������r�-����fb��J��:���g�G���0O�@��͛��.��bOOd<����Xg=����'�w��:8)\y��пM�B�;4:M$�ڴ���vp�$;c���]]}��x'��|��!J�#ǃ>!t��҂�����=8-�d�B����+ ]ez��>�u���.\�h"S����!�C��9�P!I��m閖��r�s��~Y�u��<�֣f�����	�Pq�|ɜ��/n��V�U�=�yt����b������}4c��C��.�.������ԡ�L��(�2߿+�vCVJ
\���v���Gw��mW�jy`g���Ή��GP��i�[�kxT�U�h3�H!�L��9��J��3��?'���8wz>�z�޽7�2�9��n\)�<�n��S��!sݱs�_�?�_� ��!w``���q�.��T�7��D��[*ξ�	�mu7�>�)�%�{w���H���`�+._L�� ��C�|!g[�'��N2��'y��ݿ����ͭ��>���؃tAX���Ha�0����M)ĉ�����%�}���-m8
aL$"r+IO���-[�0'�::�J�zWP�Z�5k�ق�����Y:rO9�F�@
uDH#j�3�P#bX`ú��=H���ڴ�D��Y���-�Zr���d��/����X�����S�������YK��!��1NHHׅ@+�D��T`���d^)��ƣ�/u���j��ﳜ�y�YU/��B�O���s�r��ٳgU��y[��>�=,sh	vuׅ����2.!�4aAc��r�� U�*���=1Y��'9� a?�{E�y'v��3[[JKKwg}P�Z�'=��s,�i��UK������s.)$�zY~�u�8a�X�n���H~�5e$��f3b��T�j�� 7L�����V�m�<��אg~uź�@YF8�|_��L�����@:������{��kG��f�Y��b�b0%je	k�^��Eꭍ9������P��QŴ�������ڋ�����g����Y�莬�2�(�-ح666���d68AlwMX嘛.1��� ���!�ckk����%�����8?�X���`L��!A��1�~��A���ȷkG�	 /�X.A,j0vR}=�X�,�O�n�۫&)�n�:���ܻ���\]���D"����|�]�8k@��T�����ذJoϠ�*9_R�~�E�;_?�!!�md��	֬}I� �@`�J��/���S�'q�V:��>��R7�b����.NN�7n�P �����܌��IzO胕7���V�!�{%6ԕ��W�=�� mR��pSj��/@�!�_�<
Z� �t�f�*|�0$�R� ��\ɦ��RZFF�����v��ȡt����5 �e����<�H�V$}*����c�b}�,m4mp�z��D�M/��UB���3Y�?���� �������{��*;Ҝ���4�;-llH]X?Li��7a������w3.����I���T3��q��u��*���g"aMI�ǻ�&ءz�,v���?Ӟ�h�����iƹs��f2�K�8��`�� �I�X/�y�r<��З��'i�A���i�^���{Xfa�I<-˸)UՏ��r� n�,��$�Dי�f�`9>V1&E�����%���مN�ȸ���$��/d��������226Ʒ�=����d��쬳��)$d��{_�; ���Xh�D���Ҏ�4�`�-OD��w��b�R�=�h�>�p���'����� 3&&���p�;[~)ZS�ӱ����.q�ϫ�Ӆ�42օ�b�۞����/B��YSs��e����]�<=�8��q��C�����w�ۭ_c��o֯�9>B�>���U����ps����G��.$�xA�ө�oL���U�^lJ�,�`���ަ'�΂ȓ��3��mDl(G*���q�J����R���Q��ʠ4�q��*���h2��^�`s���wW���*�Xl|�}�Aμ���d�����J�fy���3Y%y���Wa�??���a�s�H<T��*�`���މ=�K����K�3H�������q��j{>�+�#��d��С*��J8�:�"J{�[N�Ò94�9; I1����&��BAqh�W��JKWN8�b���eX�ѵ�S�x:� g���;��q����Ȇ���v�ٱu�&�+a��q�Y�T��J�kԁ�BƷoO��}�Ť�R��fł ��C~Ph;��	-F�����7or���t|SG�b�/����"m�5dk��)Dݩ���k�9T�'���cqk�#��*!ZJ��e3t�|@��E��[�=�(��4�T�CMرc��݃�� 2�|�7���E-���T~�/|��R�P��lg��3E�)&:z�3��E�lW����?�IZU>U��AC�?+k_!l�j�����R�'�.�Z>|��#����0�G������dƹ�Ϲ׻g{Br�O�y����
���:P�f��o�'�������]�'��b��\���"�Zݽ�9G��=TS[���C���:[�I,���ܼ	��W���!6k0]�!W�27x�ÁͿ�ִ���N9Ě�ۊ�({'|�ECaH�:�����,$ࣨ�Ekkk	�\�0m������	4�Vk��^_gW�D�(����c�̅q]!�O�z<�x�?���~-;��@@_��2�B0X�5���z����o�9�^\��� d��8������ �E+i���mRx�B�Ň���=7���/��>QlHc|HX���6�l�[&=�L�>C�v�gZ-�P?JnѤ~������dr�UB����n���� G���k+��xv�}T�,,,|�ZWW�����]�ڑ��N��ǟ�8;��s�κՔ����q"o�h�䓳�}������
e: E�BP��i�Xա	�r��~�@퍕����n��<'��#�W�@JJ
}���.��l�Z��H�h��E��v����	v�*믑U?Y�lŪ��㥥��9�
�*n��#B!�EP�wf��ː8�2&�!*A.N��^�1�	z8�K/�Ď�b)(F��b�� ��M�=m��F�yK�j�����-�k� ��N���x\����-;4�C,���[�d��=ˮ���pK�U�5�f��ҕ�̀�G,���.;����'dO^�{b��e�1��Re��!s�6����G��I4����<��LW�����V�=��� B���Xd}�|�Ԑ���;�����{��5����W��߃Q��KKK5	��*��פ�]�l��o>���X\[iW���܄-�������^����s<D1j3�0M�鱏#~���'~��2��^<�d�1�-n��G;B(faaa�A�*�	nS{3��,s/�A�khh���xx�b�W��1�@d�X�E?wt$�Q����1��GV����,���'�������k�m����o~�F��H�\�G����>��O��6��8�ߑ�H�3�}�nD��{�~N��[D�~5/W�Sx�5r)XChg�b�����g(ꉎ�oO��sW,�5��6/0�ӥ�X�0h�ֿУ{�3Bػ�W�2�Gw��[��P�ʟ@�=��V�ZݱL��5k �
 y/!��	�g{u�A�����'Z���ީ=Q�^X����"S33���["���wN ���Zk���E���"�������t@�Wϋ�J݈ׅn�2^�}Z,��W���t�9ͲJ��D��%���������ݻw�U�	�����tuu������
~�~����G�s�����ld_�ku��L}���o���>�g�E����633�6)��\�o�M��E�ʗVZ&l��s�I%���N":�0��"fR{f�O��La�Y_���z��D6o޼�Mz��&�N�����CO8��+����9�����Q��-q9r�)|��ʭ�g?dCqA6o�mnLa�%\V��g�r�^r)xնg�'����$H>����L�ӷ�E�#N �������EF�;����}� >����v��}���w�=��F�D��ps����(����udĘ��]*��x��Z�/�5H�aA�3r�QJ���V��X��{�h8~*�U�jY5c��=.�����<>����T�|G����U���jڋ*(pvs��X�h�����L`���!!V��Qn�QM���g�El�z ��En"���*?�1�{��4��z��D�w'�l�/#��)��R\�C����
�;!�m��yV��I��s�~&j� cdu�@��C��֫j��[<�W�'�>9�rҷ��(�7o��<���<w��	$��2 ����"������J{rrU��_��oA�d�<�r�I��F[[[^N�:T��i'["��"kb������n�Yw���P�`�[�+��&�?�{
/�����j�w��As�wt�+j~%ux�5���y��V����kv=�~w�pb	���4�g�E�똕�R�Ђ�,�~�wYt9���W��DI�TM�TU��p�p�����!<��~�H}��e�w<
�Cd1`)� �,<l��{�� � �x����BV]��0Pom��0!5Ig���ɚ����E�M$��h#S-�]0�o�z�J�h0�z��CD�C)�J�p�U�������PD�P��HF��6ke��@�̺mdg�o��h��fTYc��Ǣj�[/X��1�hWr��U�&�<�z��Z�KHHH���`$O�?�~�u7ci)��/�?V+��}(�cZ�]
hP���OC]�z�ָ1Pmt�a��Har	�6�gѦm�喋���8�ѽ�N�^��o�2���Ntf��h!��
� �/J�P�����Hm��m����j�W^��+�j �j�v�)S1#�y����U�'�ܷ��}[�) ���}�����l��i��DQ�ט���i��]�M��ˊ3�]S�5�Dc��������Onn����9�' �PO�R�V�w�� �o+E]����8�����ё6q�� x ��@|`o�W��i���n�x��<�P�>d�+��HK���̜��3�ޥ�Z������Y�!6�8(�����M�p���(��Nf'?��טzR�FGP��c�<'����S�&���Θ�4Ͱ����n���C6�Ц�QSx:��D��n�'�f��g7�K�K�$G~�N{���jdf���������^���������(m���Z�?�VTO��yE�	D��&�����l�/��%r��-~fU����O ���@Zm��w�&�T2��^8#DH�M0�[*���6��{E^AŃ���sm�:n�U^���������b����t~���C�(�3��?�M����+���%!.^��� �(��_<���O����|8'd1��:��5hb�W/Cֺ��u� ����9�R��;vm�SDj��C=�:T�n�(���A�4:a�Q�<�C���K���zj�"�l���)��y�M�/$�iCK��E�0�D�yB�����(ӷ�!����^8�EKK�(���24�>s߀��dv� �et�ֈ���ef�M:�.8��Hµ�,bN�����ߣɱdK	��P�YYA��u��g\e��JJs|�Q��#i���#�3�t�j���M������!�!����м��Z�M�i��ƹ��Ad[I�ʃ�� ̅�\ɡ��T�w>��h��R4T��ԙs]��X�4�M/+f;!��1�	�\���Ѓ��v,����E���\�֝u���Z���~[��~�*�<r�:��	����Ӆ�����6�-��p�v��`�?{�)�����߾m��%�z�u�w�����O�oX+1ao���H����ȍ��ڪ.�z�7��&c͆*>݌%��痑�/�z������h臦������Mb�!�惛'^�4�D�GT�P����+gS����A�o�$��փ~��l��4_�nUY}t4��H�UM�ު�Ws����&#��G1!��K]읱�(��x�u�f�y3�Kc��v�4����􁹹��uW�v��3����g4����sX����?8�0��~�H��L&�Ҙ�g��)�qZ� (��1�N
����=��,I���(����tx#���ӳ�	Ǿu�*YD �C���-��IYC/�MOK;P���ӿ'�TFN�f������y£��s�W����K��eOx�B��ҟU�Vꌗ����#}&p���]#RSS+g;\hR���	��&�t�cb�/�(>��ǝ:C�z ����Ü���̕{d59>�F_l�����4��B=�y��������|||^���x�E���Β��_�&��s�_/�J=�k�ܮM�1aj�r�7���'v��"�+k]S�����o�3��ծ��JTsI�~ɚ��%��r �0=��5g���^����� e�
I���R�I�'c^��s�)[B����՛�zì��MSJ������W:��9g��aUUՀ��"j������sZ��Tا��0�O���Ŧfff
	[]JiD��Ѹ�՗Q9ŢBB���4a$�Gi����Gw��]���	D�a���O79[��dg\wm�u�8��vO���̇�A��v����W/=p�m�������h~������Yb�X�5��p|����w���N��G9a�}5S��� i��e7<=��}�v�K�|NN��1�ʪ�D��`��3��۵��q8\d-ȣ@\wv&��\9�<���� {�v�L�[��Y���&&vj"�2��������0&&�	Qi�P��tгN�#8+�r��t��gyy�]��c8�|$�ʠ˝�*�ڞ�ե�$�<�� �G���$?tuu�����*���Nyy �!�yyg�H�g6?�ņYk.W`�)�°#{Y�/U��,���7�B�j�7ʊ��SS�R����#�]]��k˗ao9!>��=��DVu�}��2�<���3�&ǿV�Y٠L��f&�u�b��+2�y2|TR����dݭ��:�����~i�K5���RVR�'� �{��-Qa�Y���Y�	��Z<�;�{��0��g�q�~�����,�Aat�`���չ*`%	�9�L�+
��U ���D�T�#P��X��/t�6��V�&.9�\�����Pl>0`_l���j,�L�f�"uФ �ج5:�$�{4��8<�ٸ]�Ѯ%�n՟�p����Z�}"s�=r��������9�Ο��^x�����t�������H�~s��@�ol�(p>�6  G���Ȱ���Y<�D/��d2�<6}�����[��(�oe�`�9ͺ9�uZ8ժRC6?� YȆ�+N~�2�2���l~��i~��|��W���\&���@Y�ϓf�lbe���2�>��6Cs/��,TV����Q�.�ΙO�'Qx
��s����/�;��x�5ZV��fk1 6�E�d0�`"1��Pk�0�� ���)����X��3:xi!�����NO�@�������A��e)�U�N������+�����[ ���JP9?�+I��	G=Yݏd�kznU����������?vK��nx"ܰЏ�K�޿#R䐷��9��^��7_SI��K�V~���Ð��pU7��`]�İ���|Pĝ0�x�N�����&&�q����Se��3�HE�A:���,>5�W'�x��?��i�h_�Pd�������<�Jq;h���~폘�GA�PVV���Q�LN恐��籶9�F�b}�7�>��R����[}e���m{}݆1�*���*GQ\!�q�Hw�HYjwh�5��H�)�[�a�ҵ��u�>;�����\�&���:�#�˃Yo���z�L�>5���s�9�B
��t"�����ow�l�1B&�#ȡ�.w������@g�)+Rn��`��n�K���a"��:TK�S1�)j��x�)�:�Ͼ���c4��I�kUz唬���T�0�!��,.�*SH�-J�6�'���@�候@��ݒ2���WI�761��OL�i�,X��5�⡒?��Y��0��1�ẹ�����H�300�
L~}��9 �t&��h�/�mw-�A�E42s�&�j�$�M�{��J�|ͺ�"Qa\�)�\��"�i~�W�Gps�|��EP������ērR�>l8�x��������)��KƱa�uC
��h��&&H\�"�����ף7����f'�@�_7d������s�R�bBNr�a���-�O���]L������Ǐ�5�3�0u�w�P�n1�>�Z� �@��Q�[�$�ngJ�|K��Yʆ��P1K�x=VV|�۠��<k�֌�Ӊ��8R��  r��v�����hbz�Fg�4�3��[<k#I���[ϵL�:1"��Xу�I��Z:���ųeIN� !h��kgn��6�oO��+#+RR�=��������`��<�X�ؕ�����	��u���E]��>f�@Y�m����9�މ��yA�.|�z��[�}��.����>g'�L�g�bD�xS6q��-M􉕕��2O���ńLM�+�xA�����W �;���8��<+�Y�ҟ�T���a=�e,��~�"��P���?n:v�H:L���f��N͠�Q~y��$����G��I��Ned�, ��1��Yk@0#A�i��/���ksvr���Ҍ��F�����h��be��^]�0�:�3r��B>Vj"����V��1<`���fW~�]��T�� ��I+#���㮞�j��C����#�SGRX���b,�#�	`$�� ��r�f�e���Nj���	��MJ�{�/����㶗�<��ڂ�ܷ�ʹZJ���%~(Z����H`���$$$���#�mM�ϐ��Rԏ�\�5�����]��߲�&S'&�F�q.�����|���q�!�5�ަ��2=��#c7����qT� ;�{?).���n֝Ɛ�-�ܘG�<����w��2Z<�,����ط��H-�`Cl���5��1��3���e�Ȏ7��q�����!ͅ���v�'��l>:hLٗ�Y�OL�}�G�xғG�0Ca��1fC�B0nҐ�sԟw�7T���.�&�����x�GpۦG�w����t(��a�Y����*];u�W1�K8�+s�44�ꯇn��i=;�
+�ۯ��l�Lm`���IX<�����`j�5	����ԉ\C������&��D�z�S�Me;�%�AC��:y�*z���dc�$jT�E��yJ|���y�85�tTg-cb�.��T�&?~\�����M���)�u���b�L`j�kB^^�%��I���9T����ҳ�e�o�=Y��'�����5i���a����9aERVW�oo7_`��qݨA����(�]�>;c��k#�n19U�p�0�;����KVrv��J���~�h�Z�j�9���N�g�a�}�����Bl2��N4�Ѷ�?n�u�����8���z�#s"߰.z5�e�j�:�.��l��~��ݚ��	\��J�a����̀�Wt��S��{�|����zN�c$8\� _-|j���GO�ʙ���;L�����.P+����L=mP�;�&Qg��^+����?W`[�����M(..��AU�?��|�fG�-P��.0`��o�r~��� d��e6�>x�w^䪻�bIl�Q��|�%�e���C�(	�M72ʌa�ȁr���P�$Wy.�[�k�2E�����ى�B�|To�j���˞Rw��_��+�b�����6&-�95\��d�,�	�~{�0�;F?�I	�\^�{C��Fs�i~��G���[^�\!��摵-�1|��l��C�Ŗ%���&L��u�~�$��Ur�S�Y��-{޶�sݨ�����hV2�R
�����؃>���ц�-k����6N�����{��kHeW����&�n��
��JX6C���V��D��j���uW$�����L`YZo�'Ž�d��y�w�r����4O�JBI58��WtQZ�;�/[>f��ivb���?�h[�8�Xk���R1�pv{'�VTA�nl�4�׽�J-W� ��cc�]c({�䁫E� ��������1��Qd6B�l,�ຓ���Fjj*�{�m�:�-��uU .-�B���^>�q��
��R�o'C��B��Aڡ����3]zG$4t�õ��Cd#r���qsϡ1�k��컫כ(o�re_8�E���_�c��A�*+)�F��(L�ԫ���0�o�Qv)�i �����k�Efmnn�|�t��A���fX��n-$w�:��'��P,�e�i��������v+�LI(��{�� s��w�-�A��	!����#�]T׾YU*�Ys�� Z�?}Ux$?�������[Lo\�W�L��z�ԅ�.*��?�HD�� �~gU��e����j__�6_r� �Sq���,W����8<Z	���D�b^@�����d��T�s<���K�N�%���B�Z�W���8u�hJ}�K#I��V�\N�G�B&ygl҂SM�1�"�Q;^���l�����T�Y���0�Vn��G�-ϩ(�4BJ�
�s�կ
?�[7����Rq�Yߝk���R?~V@����1�0��v+�:�u\B��Ϝ�u�ѨP��PS&!����>����^݆�������K9���u�!MV#Θ��C\o�4��@F�!�Ԛ�L_��Dy�����=��j;��ֱ�u�4)��!�,^��� �Ӣ�:��f��� K�7��~��@�� �.�.W�=i���狭ь�AY�cv�p��&~.ed٭\�z�<|)@�H &�D��yj딇F��\��dbA�l��w$�l�z�^�b���Z��iA�e6/��N�������iC��oΎ��-F)v?O'��o1�V�SI���Ԉ�&܋�#
��j��	�:�浺��f��`�b��ߘ���V.��Z �����P��L���5�d1�$٠7���*�&'����!ӄ��.���I�Sf>Q$��V���cE�?���8���B��un�U_OOO��dc��<!$_Q�;�Hz�"67���3�0�>>>0dE})�&�Fс�*z�Z,��}[��D���э�"����a0Ôt��(�\{�Bb|��~i����X,��{�K�0�>,6(~�aܢ���:����b�;������-�r�vf�PQ��[?����g��H1�	�Y������!�3�����y;2�C�.�r�K��h����&	�K8�ŀ��Kȕ��K�`F�Q��6ZH���&��-��ie-�K���e#�1^�7
.x��ƈ.�[~������f���^��Toe�3�>Y�j��At`k<,�qB���t�٥��^��r��p����櫪��>��|ɤ����;�WZ�.������:�̍���d���NO����zK�Sb�{=��1D�2��K˱��n�/�h4L�R�z�3�9�0?�B[6�]�/r�����@�̵��9��!��;ɲ3O�},�U?��&�Ɗ�����f����B���e<=�4�������z��=��3�4�����`G��T��Q��N�ݣ4������]<Z��<��@H�[ɚ%��N։5�`��w[ͤp_�ȁ�Y�N���p�B�%�)��	��/�d�[�:Ƨ�+2=�� ���%��Γ&��8D�|%Q�y��H@3��#K˨��m^�$a�j����۷�e���j� �87a�?)!f$�* u������xc�����Z*�1�Sv�_�';OsF�N,l���S�Aff&�-�>צH�"p���e���	1����cZ�8iG��X  ?���$ѥ;Gݗ�Ks���xU���h}�n���E���$�Ђ:�z�v��~�������W�H�3��>��/8���&#���qw� 8��-_�Y/Fa�7�Td\��n����l�`��ͣ��������l.��� ߘ��Y|r_���.�4�K
F=_��X'��W�3�Q� �n"�܃%!>tQ�E�l9N���F�)�/��4���M'������x�����w��x��3G�ƀ����v����y+Z ���b��k�b<�Lt��(?�5yƗˇ����/(z&s��y �ԔӨ�@�uC��F�\�����\��%Y�$I;��?5�[K<���Q��a)}����~E���}\{��=uMp���^|����-�h#u���6���q�K�Tu�{#�dJ=?a#M�4�\�&�9����O�0�܇�۹�c��Ų��R	��.ץ|�6���AP%*>OL����b�sK
��ƹJ��v��ɽ��!Gre<�vC^�����Tb��h������\|�J��H%y����j$6�Y�v���4���'j�[��` 3u��4===��F���[�+#��Ej"3�Q$U��2`$��EB�U3�ѿf[J_��m�)���eaˆ�/��fX�=�HM�0k,W�L,@6�)¿0a��Ś��9a,�z���cf�ឣ�^I�',;@-������"�A���k+
�k�`3N��IAUY
�[�\,��Q��/)V4(�ߴ�fi۞�[���
�j�Z�w��{�^��~�� ���¹��k:�`�n��9|���o�y���Ԩ�G��|��0����K��O�D�����1�P�C���H�+�T>�jE
��UM��i*�5�S�l�3\�����b����'c��!�v9�Z�A�!� ;���'������/��Ҋ�1u&]Ⱦ��Hx&�ekE��S�͞?.
ױ�	�S�� �r��~�c��C��8p��:~��P��vlk��W�����|Þ���{i���>{~f0��u�s?-��B���ϼ7���5h��@u�[`U�D��Ba2(�}�
�-�\��9SD�3CS��%�w6�t�,O�P5��s���J�{7���ŗd�}�<�� ��g��Z�Ref3�Ni���R����U�.��ʣu�8d�XzGuW w!��|��ʔ|�D4��s��!�p�N��]�;�w�k�0	�cMw�_������͈ل�O����;�����3)�qj��zH(�w�p:��ڱ���~%�r���Nmc�Rt�bL0��}�^#݃��[h�:s�'?�ԟ<��0��/>��Z�3��A)��
x ���{���y9�D.�;�X��E7߃�~��m�"Yu�q%���w�?��2]�7z��|ȏY����0�J��9���:T����s���	%���u�%&�f��I7�qO]5n�3;F'��4ߤ�w"<�k~�]kjh��}��c��G�R�p_�:E��}�����-��-\��O�x$��zc6t��#��wgR��H�Xk�F��}�0SFhEڬ�˞Ho��~�$<�L��+A�Jc�i~z�3�e�1l+��yz��Y�d"��rZ�2�1�D�z�^w�V�K����_�t� 9��1���v>�g��CC�@j��� �p3��Φ97g�:C�;�X�&��R1H	�Jk�zr���+��@����G����R������ y.eV���֟|���?��}�g/�j�m��]?���d0Fal�c��e�P#���2�vy�����v�lj�"�D8��BN$��0���l:��x�𽷊����ja�\X�|��~5��A�%��C��A�W�p��I1I��%��-�sy(J9�r ���HpB�b�K��M�[��'�ո���dwL-�ֲe�ز�];u_�*h�!�)��M~�֐tġ���+0j�U��kE��q��.��c��#�_��twu���ƸI�;��	�j*
�Θ3d�ko�Z�IZ�h!�n�H.,�Mj_o
�T�����5H��
��w{�-pq�5��o8z���_Q� �����>�x*�A�l��$��i*@ق�r�1Y�;1w0Q�j!2C!um��e���R���Y/�fd�
�Wm.�h�h���V�H��� �O��a�������TG���@X���WF\s�WL hN�G})H#��W1Z;���j|��R����)��k�JY@�7��K��pb�|;g t�9�L3�/W��g����i�Ɍk�-�9��;"Q��6��M���?3d?[0�b�0��
���`����&<O<N�ӁQ�%AĹYw���V���y6G��z'���v�hf�$Cf���l����_�����I(���g���HOҗ��3����� �����=חH�bm/i�>=yTW��p��J=��;�?8W��V��c�wq*���m��[;�Ԓ�!�)�FWA����C8���\oL�v�r��s��u*F|�=�e�8�ɮ��5�IԏQ�7#_^x��B�P�HL�#�틘fÅ6AG�<}����l� �+�����QYj3�����>�v^ߩ�ły1m8�F��Pl>;;{���	巻& ���	���X��
y~���I9�B#���bS*5��:$�p��H"���F��������ݱ���B�.͋{@}����亦�Pz#$�B��H��'ǔ�֎�?��V�.��=����]�x�(�ȴp�h��5��Y
�p1�7O�[DXxs%����9XÐ䓢ƒ�M��ߐ��3̓ѐ��Q��l�ch�}�e*�\C(
)n��a�1QL�n�d�+�`c:!��<��n�L��9��ׯ�ӻ�����	�~���&��#J�&�o/z���A"�"��ul�'cWLmJp 3],��*}D:޳�[Ik����]j����{�.��F&�=���Mf�v��vx'��)�SV���J���F�.�sM��f��0M�p2�l���p��D��]��e�:3��(ٙf���Da:7��;iQ����ِ��(��P��=K�`Z�,Q�����/���፵j���П���7�l�l�}1���ۑZ����g(��w�t����p�H��>v	

��%�£h4k�맹�N��#��#Ғ�� ��9f�X_	��`�Rwi�U�9����)mo)s51����D�&e��e��̗���U�Z\La����mq~�,n�Z�{��6�n�ǹ�[���ϙ߸�ȝ��� �n]˽����SnO���> �o�]���]���]���]���]���]���]�_�|�6������$*	=؁qA�ڽ�ՃE����S��}�(����}�鍸 �5>]O<��^9�X׷�r�Ӵ"���S�CgB�>.?\饪w��N��3T�͒OoM�%��A]/x!V����EmE������n���o�o[Ł����ԼZDD�,��� !,��c��!��%ߌЃnTgt�\l접�bB��*!ʾ�jj��?�;ܘm�����=�.FvL�O�>=7c$5����Cʣ��&������4Fy�0���q�����za�3��ɰv�Ԡ
uji�~�W�ƴ���ٞ@�y������kI٩z����T��6r��_��G��<�/�D�+�Z~����]�]�OClC�go���?}O�.��L�~6h[��ݒ4÷��Eb��ٱ�'?���E�/�ut���5����c��u?ߔGƞړ�޽{��UR���
]?U�PK`:&.Hs�~Xj��9B����@�����3�����x�Y\��]�������~��av�ҋ����&�7:z�h��߼<U΋���y���x��b�޵�\X����KW����3qu��UT򚚚���������(�bm
���n�õ��C����277��pUEⰒң��K����+�z�߃JZ-Je˖,��[R��e�E�˾d�-WFH��k��%	I�-�l1!ː��s����<���^w�|��,��}�9�s��Ae���P	q�"�Sm'�Dp׋0Aѷ�d0��V������o��AwL�C�S��?ݽ�\�2rKȤTĭE�:����A����OOO�\���b���H>��l�o߿��GO[������0�KPRR�-�ū^�RB�Zf�R���u=	�7�m"''w&if�/k�� ǈCǴ����zk>~������gҳI��A_�p�ب�Ěw��.G�����߭<+�u�����/�^�#���>�%����=������0e�9vqЏ2m�=c�NZ�5�r8@�����P�
�ء-�d0�\�GOO�R������~mӊ.���[ξ�fX[ض��J\������f-�D���� ���x�b��EN��G�^�4u�������$����<UO;�'<�70J���X{��s��vN����uҹ�
ї[H�~�ܑ詟��e�%�`�}u5��{O֩Li���*�[{K6�q��4U�W�C����*�����W��OSjB,M�[�����6*A������ס_9��)V�R�s*��ކuuu�5�5&B1Ȩ�%���Mۋ�0�4��)�K��9t��ԔQߌS	�#�f"�oF�������9���"�Z��_�1�7�S��ÿG�r3���{z�0pȦߦ�˯�x����՟��Ԥd��1ͦ\�>�[l��ۅ._IҼ~��QLLڭ[�b��s�;��<���Os�;K ���W���'?%��mZ9:�����Ν3%C��}łvN�02;Kij��!:W�4�ɹ!!!LE%�㏻	��=-�G����34�a�`7u9;�Y1�Y���-J���C�FvtD�hK�zt����e�r��a�
�9}����EuJ�9%����af�/���)��ߍ�������?_=���6^Pݘ���'�^���]����n�O\+د��s�<���+�y��G>������s�P���TEԇ��#�`\�ͮe���׻�SVj6� �Sl�̞]�|�Z #2��o_#<%"�Ã���p],��m*/��o�'�c�dÙ�
GG��ч2��^镕��϶xj�@��(����KН�8��3��TxC�NݺS�RP�{�M܄�<:Č������{�><:�d����!'���zq���L�˶~*��  ���"�ɰ "}�'Ff���|FFƜ�1Ew���ulm3.����֏������c-�̳�ۄ��^�PZ�?�x@�?�xb��]�\�KE�K�_D'��Ss(O�'U�_����2�?�IO���x=�������	U|a���#�vU��~;���o��;���f�����Ь 
Q��ݯ4�T�M�1��k��S�~�C���n�W91�)]䁮�Y�۷����`VT�O��1�r�-6 }�Q���R��,��2��1ְi+�}^U*�H��C�/^����g�G��t�;RK�%jh.�u��ۊE���*���C��o��ej�����",Gp�O=����7*�xT���xt�!�z����͹2i~�F�S&<f||�_Pp�����M^���%W�Ʌ]]�>�	��D_G,@�2�n��[���jd�E���q�/�6EP��X��:��^�3��Z2$H�UoP[�q���; "�����g�͍�2��� D��_�;���}�SQy��f8t�&��m:R��c*�f-E���u��|]Tx�KCA����!' �jk����MP������ڈ�u�o��l����|������U��Tk�+���8;
�H��\��^�s��1�YL��/��~�J�@DWb��׍���ff�k�1���]��y��mtf&77�	,#�������ʢ/!���)efh=g������u[������2��.�<���h����ľ�)���r���N@-t��w�P�X�|�����9�n�\Zm43'�v�jiY�c�(8E��� �y��`�ݡu��Vp��Z�����"�W�nQ#�cߕ�u�@��NY9Z=M�pc��vt�%X��dP�B8`����-Kkv����;<��ia���o��r��1��@Wt��s���[G|�N!߳9�ξ�<ۙ�"\'-�'T!� xu �m�v��$�hyʔ�0Q4詈��n3?5ڽ�����7n�*�gj���y��ׅ�Nx��hu���k�sKE
�.g�XB�Ɡn|s9�U�g`+���.����a�� ���ƅ	��Ww�m}���'15tW`^��}�X�}(kk7;;:ҫ�QR�K���n\;�:�F���������/�սx썅frrrܓ'�ַ�&Z�Ey�j���4W�S�������þ����/D��.�Qd ����|ɣa�-r��v��Ma�r���@̽�7Z-�7��yV毙㓼��|1�'�Sҗ�-3�=��x�����\C��߷��G_6�V`����l�9/�b�?���swͺ$
V�mK:��@(� !!�g���J"�����<�"����2Z����ILX[z���`#�`���j�>|��@4Ǽ���e��3�K+����	ɚ�>��FI����"�6/��oss�h�Wq8�xˢt���<�VN��@`�u�������f�#bbx`��>�P%�F�[�0�zu���ΐ��C��$%xfT̖�X[[㺶p���S�@\V��ֱNDWG'���>Uf*��m�\��!��[=�#.P����]��kij�x�cܹ�chȹ9cž;�S�fU�2n�~�/��˪.ʹWn�`Ƃ޼��jm��=�oz��DRaz
^&1V=��rp=2��[�<�v!�t8̼��1��n{r�}h]Ry�4����E[`��f�^��萙�L�9���^�:��][�nr���<���ﯧgf�
=�^@�u����4[��d]�Ƃ�Ү"�����M�^y�cv|r��Q8/?�?�sK~aa�2@���坌v���i�[��p�}�.��N�XM�j3c\�z\w��a�`:::�:���������tM��m�gb?�>��*��@�So��{�n5Ё/+e�+Qw�>��·���ʁ�������-���K�~���9�)N+�-{j�l���I���U����*&FF���[޲������4��@�-'�t��Y�fyKƕ�jE/(H&��֛�������f�h�8% �!����D����<o;��Fƌ�\�X�;1.N��U�,���(B��`�-���2��I��y�ec��ⱸ���#Q���!�&�(a��vaqQ4������z�G�~�omj G;�\6�D�+P"�rM�mM�v� ��޽υ�U�;���W�;��O�)�K��)|������5��X�#.� ��XD0���ã �`PX�?u�ĕ{W���rTהn4�㺶���#����^y�>�챩�F F���^��~��!N|�k���!�p+��tu�ZFF��tu55-T�D3�>6󔳅$�L�\������?����(kgi����~��~)9b�(��B�K�����\U��������\��Fط�0�����ۨq]Ŏ��D�聦-�w���<���'GA�gܥ;{z�SS���7O_�YZg���*d�ˇqW�i���*\wx�(R�>�M��4˫^'��!�����L�2oq����Ϲ�ПF�ݣ�H\GGw�����"XYi�n�u-�ބL-p�*�Ou�o�	�!,&��g{0v��j���3��!Q
�C,ӓ��X҃\��H;7D0I�&�˭b���)HcY���tP��+d�Rs�<g��w8#���R _J2J��Չx\�6��]ۖ8 m�l�j:@|���]\ǻ�S�JJw@L	�跈�A��H�8<�{�T�c���G)�-3}���Kc���͸.AQ� �wݨ���m��}v��A�rsZ�s�46^����J��|���f�++�@���Գ���PQ��~�����������E#}����AVJJ}A� 8;t�`) �E.����qܔ����?4X�d�;1q�B�٨0�b��lw��mW�|@!���o1�G-+3���h���"���,!I/^p��;�	O��51��v��zZ5�3o:�b�@,j���ڧ�&X߯�xН�*&ff{ �����Owi���K�Ʒ�mx��L�\��%�)',��������`�龜��3SSm^Ջ���,�N��:^����[��u��a�������%٩q V�J�X�>�ڗ���� ��@L�xdxi��`KT����}}}��^k<Z�ʝl`棄n�,��8:�N��Sc�?�u�	��o��n>������������6��ي9y�#��)w��r��B��~���&+Q虁�F8�_�(��wW.��RПEc�F�2j�bT�砏P�W��M���,�]�X�cg�k��r�G�=��錴B�'Z�/���Y��i�`v~���#�'��`FJ\���|vv��Jȩ�f��t~�6��G���DX:�΅�-�v~:�( �Z�ā��N�T����3%s��J�f��3�
(�2h^C�qFt#kl���-��̜N5������z���1�S��rZMU�:t�*C!�ʓ�z��ǂ�HWt5𾢒���n�2�Dg�i�R#O��>�EJ���Ci�K�m���e��։�P�ah�ro��r������u�f\����>7�SAy�����??`�� E��[�$m �i80�A�|�����;ڝ�?�����%�]cc�s�N%�}}H���Q��KӐ<�^Y�!�9UL�m�\=����QVP�dm�"���C�G�764��>���}ud:���̬,=-�羰B�C�P2�~�����D���\SRV����;�Ae!~���Z_t���:�����*��}Ŏ:��S��}�}�x���<�����{�����$i�<������8v��K��A�ij����Т������A�f���q4L�ʉ��\�_�.�32b	�����bj�]��8�4��w�V� z�����b+�sl[��@��9:�yxY{P� +�D�W�e��j��`��� B�u;:V���&����a<Y&��v�O��h~�-DA�Ģ()�����eTV�?���d�%�ŏg|'bm�.���3}%Y/��D� J�u����Z46��|(ӐH�R�ulA1(��н� ^�N�gA3mϾP�g���r~ˆ҇���5gff2��+�^�{���а9R�t�@��gt���9dl��w������'C(q��<3'g&D�Ԗ1�$���A��
dٲ�����}�ƺ�r�g�No�<9��w�m�$�Nw��K� 4���{�ߥ���J%//{223c���wSy��S�fa���'<�ݿ!����َ5�|ǁrbȭ`��oߞ��3��(q05��[��X޽gOYx7�X�)fţ�q_��\��}%���g@� l��{�I�+5�5C@L����f����o7��BPfTT`�Z�LDCd�����:��a�9!fd�����@��_�t��lȀ��&�T��ۂqK�;��#\�������;u�������-���I�%mmZ��e��N���v�����������V:�}�LU��ւ�Ru��7��Ԡ����3�a�*%` p��;&)@��?���RRlM�CVEE_{���q�4���MHA�k��y��F�����v*�V��n��k�m�m�٫i���'�JO�2Tݫ��?�=J���e���wͣ�,�E�z!c�yx6��//�j\+���]*]���DHx�XU;�Vw���W����g�\5��S����5���D��K�uE �T n�q�a�D|t7�*����R�o�e>�0��TP3H�B �{�-䒌 y������4�y%%2^�)*19X,6
���F����tHH����]Y:�z���y=��Mx� )����e��v�h�7Mtp=�M�w�V�gpJڇ�'�*5H�n���9�Y1�.$�/ !B��R�J���4�j$���{�>'��뺹�>)̦���������<��Fju"��/p8���..�����H��[���7�AYlq�6JW�	��������>�V�j���z���V�
�I��v������q��||m�3}@E�M9�����L���bd��A���Y`���e?�Yii=jjjBO��:�2}{�<��n�������[��-�	�BLM��@�`��Y�2`�qq��Ӏ{ cs�?�`�����5��h�2�l�[�.{�O9���AAA\ǖM�km���3[6ɑ ��-,,��-,,0������c�~=B�.~�\l�r7��+�ˁ�PJ�R�`�6=ݎ��q��4�ǆ�(���Ye��}��Gd%+�w�v�!���?�}U!=ݏ�!J�-�wn��+)��WS%d��^
�ۑ|��=oԭ�t:�Z\𲷲zWby�.�8یG���m����������t@���,���(�g�Tf(O�<���rGo�� �Xp���)�����/�A�֕�����Wa"�}K�����#.=�E�%���?f-��R�u���>d�_jS.�,��{VnU_Ymhn��j8ߣ��(�l Ef?^�m�KK��/]����˶������ܹ����%K��	ʱɫ�繒��� � �!��h�U4���a),tc���2�R�������u� fɱmx1��� �+��@c(��ڟ�]�G<�K�A�l����V���(Kxߑ;�hJ��T(�ر/���}{���#�hJ���!��!�W���,�3�����J���oƺm\o��#!�ϻ%��V*��FB9��(f�Z���֕g^�\1�D�� �|�v3��C�=	,c�tX-ԁ��SP�j�
<�s�G7�:::7.��3�lw�a
?��u���t�I~�ϋ�@ׯ�	�p)Cw�\�bŷ
�:���i4\����S�L�����7�m�I~)���P��$AQپ��mhh����Hc�����wL?Ozݸ�
�#�A�2T��de=����]��[����T<�ܴ�]��[�>d�AK��'��z"-#uW���"e
?{��? ����x�"�͡U(A�T����������6�C[XE8�X�R2�TQ����ܺM,6�Ύi9�h�10�s��.�n���׮�|i���+#Sfz����EH㕡@�T�TR\�{2���_ܴ���]����{�ǧ��x�������SSZ�	���A�����Ɵ�b�S��߽zS^E����{���v�O�$>�&e�HC��F�� ��a�~C�gh&I� ���8X��_y�S�)*h-#�Ɛ�,���B�)~�B����_��H�BҞ�6����E
��
���A�gfj���oqc�S3 b�6��(�25��H� D+�@�Mjk����_�Ʒ�c"PQ�<g���44���732*{>�/�(d^�}��rJ:�>J=����ֶ]�0؇OX�����P�y�����Z���t߀�\TH�cnn�DK<�!'��r���7�S�1L��q���ݒ�-�Z;Tm�����=�o�7��E"䙱13��0����J�� ��������IOI�^<Q\M�K*~�;{������oz�����K� �_=O��m�(&�ދ���D1.� ���7��hq����4��!��Qd"�l���o���`�Rs)3�-v�G���}�_H;c����������j��\f^^k{9~d����^>^=�cu��9�B���vԘ;p7�ʲ`�X �܏Z���-��<��;���߇��9�20`�q��^��=�G�[Z[K�����sXԋ��h����P{9��d�xbX�(rDjj��)M�J�B+��IvW/�\�����Ȟ���>`�M����_	�НW3�j�YRҽ��Ъ��Uo��,., ��_e���v�
��k{�ɹZ����
C(v��a����k&^����_�ӿ�ʝ�y�f��<�r�p3�p��9NDs�(m�L��x�R��Q5k�v��c��
�;��*d�2Й��]\~ĵ�k�
���QX���߫���3X�O}���UC6m6JW�9U-ĂO���랬���۷o≈Q��L��������>�����?�>����,_���̬�y�w�%��Fm�;��s�~M���,�������{�8ǥ>��pif�f%�)��Z�������@[��L�v��a�55C1�e,��M�5;�H�\���!����=[��<��HƂ2w�u����� S����Vﰐڹ�z�۷�	��oa�8��S�U\)�n��=��� � ƫ��=�Ɩ���%(~����e�����ZW4}������{Z��g��[�ܚҟ�݂�j�iz��J�=ܿ_����湴�4@��9M����Z`��8�=�
� �m+ﯻ��4���(�DN�NBZ$X�v�:e��P9}�5-M����?����nnVZC��j?	�������rPx�kB#Obae.�?�ZGf)7�~����j��zwJ�i���F���V�Y ��̯v7�� .}�"����Y�N.ڢj��YR驧�!��F���x�<�<�⒒Y��]���g�[�����Ӕ�4��	�����t͵����	���]��UX�f4CV-�\��UT\l��-�[r���{YTbm��;�H��{�Bo}}=�y�W�$������Rn�V���@���R	����v�fr�������y��싅|D@�����/B��� `]	�u���
��C��.
�f��WY�P�޿��L�=�A��,�G�y���&(�����"9��b�/\�g�Π=w���'��T�o���l�q8$	M:>^��>W�Q��(��'j�Ѳ���s�t��5UM��y��@�W�,R.��!�?wtt�%�;9!�/H���/��F�����Z��Z���YY��>>>����V*[UC��-�A
�O��4���VbA�����������<����B�=�=�����E�h����ۜ�֦EOOo4�f�!�/�k^�)Q�sl�N�P��)���$�D
ư���*�C#`�`�B��B/~Hַj0ky���ʉc��pG�I'<[��u��R�[G+E�4�[J����M4CR$���,wbb"K���Ȉe�ͩ��U�к$P��;'àҗO>�C��.��fn�
M�����������:��@�`!��t����5Z��$�N�%���׻��D
��͖)�'�.�r�+C�Y�,ʟ��j�v}�[5�?����O{|�����pׇ��A��"��t��_a4��՘��3b�b��3RR�ɀ ���p�v�w��%9H�̝A�M�W�U��ds���G��l�΂�F�%���_/^'*ބ����Ń�v����1+Q�S�9L^�����')���N��w}n~��8I\L��ǡQA\H��
Ph�����^�B򉪹� #���8�,��z�bT<��A�o�en���7���LVq���UB�p��0�,�30�k����A3��鞨��� {�ݥ}��j���-䏐v�t�U��B�a`.���
�TT�1wi���r�%555��r�x \�.9t���� j�m4Ui@��6lQ][�Y�!�s�FV^u&��ҧ͆��E�S<C҅d�f{�,עq�Od�S�gTl�W�?��j����K�0���
�L�t��-�P0�8���stLX	����g������"d�����:��T�5�u� ����a��i֢��o����������NR�1�/��da��~5��˙:ۜ�O�ӈ�_��n݂J��K�î'2G���E���K��"��h8�V�	5�H$���d��}�"V�*."b���? �"53����������G�S؅<�I�=X�in��/,�Z1P�0m�Vڰ[�O����9|������Q��r������`�I�܊���� :*?�K���f��sC�k�+�QW�ڒ�]�����>�гM�7����:����Yۏny�0Y�V\,�%ťfpR�)����� ��O�@�ܦ��3��������
R$��������b�O+T��Ҷ�cA�Ν�]jSv���dC�RTG�Z�$���̂�O~`<���i�b"�H	��Y�����������!� � �ߋ��Qd}����0��i``��+@ϠL׉8LQ@'|��Y,��ݽ��j��u�LZ���% ����ɪ!<�*�Ӎ�%����Gp8�_[��_�.��R�G0	�G�à��H�t�}���&5������S-��оڦ���ؗ���grhӶ#�j��>�����#.h^=��������]��#�����m�"��3��kg�>�����0\���HS������OVy��SaIԆ���9���YT���{���͉qځb<%Ƭ=C'�!����#5�	�����?Y4��Lbecs$Ty͙���7w����'��>��_�<����t�^yE��)�a��������'?�2�]���B�Ho�<؂�,�B��x��,�\�]�����)�J�F�*�6U��1ƕ;����WT��c����r�R��n��Ο� (Q�w�PЦH))��*䋎������s�r+O�/. _�:_�j�v����K�|�W�1��>b�
�qb�$Fw.^± gel�e����/[�\��F���z.&��顗K��;��XE�_����붶��ǡ�j����O�4M-���g�+s�g��#1+3�t�Y�t�/M�T��e��n�����@�:V��ˤ��oYbՏ�IGY�
G����6�'�����(E8(>��z/
&�, �:.>ޚ%D�Jߑ.ߴ�#u
�I/�!v��=�$�/�����"��Q��,�TU?��vX]]-&|���0��,<@�#��H�Ñ����_�'G���27Ot��2<���u�O~���"KrJZ'G_�m>[\Jʖ,y���ޖ�����䱃��1��ƴ��9����?.���c�U3��i��bT�̜��E3x�vF8��arವ܉%R~ܥ��|s���6�!G��߅6�
@�j�\*vo^w�v)�&	_�:$vP��ħ��N���Ҟ�Avvvߩ���?��-�	Pۀ2:� ԉ\3M|�$��NC I���/��sE(���0�_���k�!yD�I!���=�f�����=T�#����o��+*��Dk[h�����ݧ4��ۡ�f[��bç��P�-v������F�	v��k-�eN}�<v����!z����w}u�qF�cSS�QwS���D�smm��V��k#�����-��w#A[�������0N��2PT�T�/���7���k3@���&$��1AY�ĴŦf$�������C<N~�듙���iV�x�����;U�f�T�D$�U�/_���s�[Ip�Փ�*��zu���.by�4B�^2�}����9��<��@9��ě�r䦧�ǈ�6�I���T�OyN�8�KH����8���`��3j:�
��S��r #�F>=xo�]��"jn����ts{MW���%����Gmx =��f(��o������9D���4m>��{!�k��>y�)ƚ�Q��q�W��X�����?���ӝ���g^9HKy}�j�?���\�avW���\�cb�z�h�9�\(�2���ə;���T� �����E@�^�~?��+__I�p$�h�F��y�g��,G8�]p��!�L��k�E��ꑮ7}�97(��j���ŗX�e�c������dVR�e���ҝ:K����yo����׹}r�������%���E1��X�ll��~~4~&8�XzMM`������٩�@)op��
tIJC� �m�l%ZYIu��۷���1v��}���O,=0_{۵eO<.�.t/�+��+ ���A�&�u��D��w���A\�M �Q���7WeC�����Aν/��a@9p�u�^zz�����Mn�ޯz�\'���n�{��.?�i���U���ZP%�rFL�^,�T_W�ef&����X�����L�����}	�}d1		��z�8H��AԶ�K��8K�	i�*�g�p�6_��x?��*lT�s��9��..5$$�af�����K@Zʫ5��,������`
�S+F=�qXY�k��u��������o�m)R)�����7{��U�S�qK�]�;M�6/�j5���ps
op����
{���I������ߜ?y�����ey芠���
��mZ{���x70ٳ���y��l�n���k,!���s�va ���?ѫ8��fh0N+���I (�{�p�=�D��`��H` (̽ T ���zތ�S��쩙_K�=`W�f�}��c7��8������?�����>�4�/^�lb�`ge-�3�{��'%@)��T.�f dy--�$޼�ǉ�bvV�Fc>ie��w2����h~�p�>?�пk]s2`�̬��U+#u��Z-����Zv2�Q�	S[�|8�j�0Gt��WyWGG!o챩e�U�lu��.������'�Ur�-v�#['�ޤ$%�Y�N�]��c���۬3�h�.&�W��_m�j����(u�/�7#S�`(�н��U{�:�Q����i�P&���c�M�ITMh��ɢ�,Zd�ZIQ�Y����ՏN;C��Ҙ�ܨ��k����f��KK��װ���=�9in��0��}O��9���.��BOf	9m����g�L�X��Q��~W���X
X�b��)��RCP
��T/k�^y��P�=����}Pk�6�R,iؑ���>���,p}Ui���, ��G�-�0��Ra�˗/C�q�������iX�RWq�G�}&��T�V��aj�sWɋ����~����;���5��T�$��##�U�ي�Y�'!��d�}Tk��7���g��mȤ���ڮ_`������]�����)������#w5{��3��}o�/~����{��{,`w[d�R�����q�ǒ���H��6�w��%/��犖[N�3����>@���O9�gC؜x�g(x���&�MO�n��PJ؝q�{<xp���$ǡ�A�%�*v�~�Y���ʟ�%�_�0-���36��u�m�7����P�������Hh��h<�_^%��=�6�?=�:8���k�s�hXJJ�7�Q#�׿̲��^���z�Md��Kn�&�������U�������g>��̣����9��e�LLL
���z͚���t���<2�䵸���n�7B�����S�7W:����[/�p�8��Bǆ��oWcH���|��U��}3������νa�9����1��C���Չ&���ש%4�����V�Z���%�����4�M|���\Rc�d��>55�Қ����ݭbĖ�;c�Ɂ|s~�U����Z"�٤�X�o)��ײ�gj(}5��9_�|9��mb��WxfJ6�nk{�6ݎ�-�����;�R��7�afy���o] �Β�~�{4�O>Q�#3�#xz�]�ЋU��n2k�2^'ńu�nߒ��Yo\NQu�[:[Nx1�>�챾��8���)��m{t�� �����L����-)�t���<"�{q�BD��a�s`�N��e�z�w�S>{*b�0�IQ�y��3����슌eԙ��|ك$��y�{Jȭ�-,��s~w]��Q���,6n�؛��Y�jU3�[�M~�.ذ�tBK+�^���iwq��oqxUD�q����^.jwz��u����D}�}3(HM��x?%Ȕ����$�0Qf�T�6�{N�:5oH4H�)��{�.<8Lt`g*�i�,1�3�z�J��Wџ������G������.��=��OL2�<M+�ߘWP����d�?��!gZ�w_�~��t��T�-+d�����]9{�) ]�R\�0�.=?�X��E�j��Yma�ۑ��	����j|"�����F�_e���Lkb�8���1� �x�R����ڸ���-�T6���+�^�u����!�ܹ�޵�����v!%��#�K�o��/�o�&�� GRA�~ҿ��[;�[�����
�
�L0���d~��Uua����`S{{�6�2�-����6��l	��;`�f`J9d��}C�;J��&�F�`b�@���K"�5�v�p��%y��]��-�XU__�e�v����1��ͫ�-o�;��6�.f�� 0a�#O�t��u�U��X[���h�.�#OD5x���#i���Tt=l�+^���5k��G��R�a����h���<첷ظ�,�C,��>�A���0�����v�v�S����Rm������UKˤ�"N��knRo�*���l�K�y�(����s��f�x���4�z.A�
��`�2�G��Eq��o�vuu]6�Lw*a#�%��k�w���E������gu<f�Aa��-AMCÙS��\;^�Sp�z�8W5h���36�M����5\� �%��6gT�D[���Feaᘻ��^�`��yӏo�Ὓ�v>���{��8g�7SO����@�V,���%�W~x�^FFF{������cfڔ9�@p��������UEE±g�D�.������Ӻk��[�f@\;{���p9��8潘m������+��H���A$`���lvt��/�ޏ޸9)3������q��Ys�zZ1�t8��#���3�~}��DeIߒSr7y�Iug�����eS7�7��w���B��D�k�������"5p�ܚ{!��W�Wj8mZ�	z�I:���'��5Rr)Us�ί-6�il
�w�t�e[ll�ݻ����o,4�I�r�3�G�|Ōs�31U1��� ����9]ōM�3#3��/x��.'˳�]�>��]�)�iF9�n���[�x|`W8f�rI_����{��9-#��&�h.q�/[���B+������)�R�����Cr��OE��k�'�]_�����״���4��>Vn�Ft�m��V�E�7~������6sw�&���H:��{� ��}��ț���H*���˗��k�(�6j@��n���y���Q����*���uE�%�z��3�f�?����־���3T��ᗽ$^b�) _s莗�D�l��y�t-��B#�
�ے���ծ���t���y� �ے���'ܷy擺ES,�����rF��Kۅ�!�m���9gzI��Clll�_Q<�Wg�j���ӛ�.�<0P=���u�]��r���a���Sp��1]���Z�Кڔ���Z��۴�߶����Zt�)G?����W�����"�Y�������z�
cQ3��%�)j$�}�בz�5��5� �H��(�N(�����������Bss3x֩$��V*i���U��<CԦ����������xR��i�˱g����홗ް{� ��$Mg��ɔ���υpǜ�z�z������Z�`��|���L���!š��!���u(޹L�4F���c�.ԗ�ڈ}�ė ���W�d�����([�_�zs�_�)8l.p���WQZʲ����nhb�~����������{6����� ��n������h�c?SP#m3��\�K>��� S���S�[Z�;:t�y���t4����D ^�oi
ۧ���<�f<���i�[g�6c�J՜��&9:���S�_ꢍK�&�[���ϊ�>�Ȯ�_S��4�Rc5 4�Ibb�^H������}3�2P'T������	~�A�j�Ο\�s�h!D�R=#e�S<�?�7�OU�aF�R�54��2&�7l�׼ߡӟxs��a3��#� ��^XH��!�2����qo_ѥ�Q�sJ#0����������C��?��S�5�j�G�$�?��y���H;�0�@U5�Ø�Q�D1"��V��	i��P	��5���Bϡ���B�5k�7�;2N�����֋�S�@��R��{�>�8_�����Σ?��>D/����79�^�&��x��Q��ov����ѱ��K]f0����;z���ޑH���<�J@��~
#c�VM�.$����jl����6�rU���NÃ:U�Y�n�%�[>}��U�b�T�N������,��!�5���%�������]���v�'���<�^UXK���j5��� �ba}v�:%n�@�z|��'Q�X"Ba�����`jj�k׸��
��@Cw�Z�D��,�/�7d����(���/�����V>�������T�޷"�� g�^����9������3��7!�����9
��6����5���gm�@�=�_��_�L%R��4v�#ú��F�v� �ɚ�Hm�s6�A�-�q��|������1G#Χ�/�����fo@���Qs�
�V�E��`N�C�4.Ҵ�Rr������l�R�Yl./,�5x�}l��Q�	�&䣚δ�F��X���T���É��A��U+ğ��?C�6�0Q�Y"S��W'#sc�c�"����w�ȸQ�%ǻ�c*��ǈ������"������Γ�7���#���"�~�x>�[gv��o�ҍ{f!��7d���!/$k��Kg �k�4⨮炔�z�Ib�"He�?�;5�(
�\�b@{\|۾�0����VN��mtp�p�+�0f�X�F�B$Kxå�#�R���54 7.�����(i����R�a��v7q���N�7�3�	'��ܿ�3���mvd:����F���bu��km)�ڜ�/�"I����:�JUA��<"�n����EE����Kg>~��Ms�H��m_�IS�R�N�����[Zb�Z���kn%���)b�f���-���w����^���h��J�³j[
�e�vG$ԏKgd7�/u�� i��/6:�w=+r�Ntέ$����-��VƈF�P �����#�s�攳:/Ǎt�q�F�Zy4� m�{����{�X�B����U�G9!�R�8��A����Lx�FoT.������J����B`v�~SF�$�2�0�
�����>�N�iص'淹�;�?�=<�$��/%�8�^�5���p�l�!��N��"i�)"��[(�R�F����1<0�p�I�#�!F�D�s��j[q�U��l@��U�S���e}���zT=��x��R�W&
i��l��d�c!��l��H��ٽ7�
�����n|�QPa���m^A�M��~s,�K�>d�E��G.�QُC�&����h��Q�.{ǎ�����z�x~�#xx�EGY����� �iϊ�����\\@#"�͖�>8ȸ�������<�����}1�j�5��C��،��`�X��v��Qڲ�J`X!�����{����T*R�m�I*7�iT����鷟>����'7���ݒٷ��Ș�e֣1l�&�6[�;u#�!�s��n��)�灆EGG�����~���Kx�o��6N��ߒ��mBڿ�g�M��T�_:>>��3V�Y�i�*4kԱ_b\�r
����m?T����;��L�@j��!26]�2�E���O�Q�B�8b<��vl�J�|A�u�՗{�X�u���:�rG�{ն��*��c�&�H���ze\uh�q����/������06b�1}����<�3��8S�p[�mx00���D� 0���E��;���\��bbt�7�KSs�Xl�ۥ��?\���� MM��-����&9���.�m�
�i��/���҃+����Prl������NE�ݳ�]~W�i���`�fGN���]*�%�Ner1���J�xK�X/�{���t��q�g���g�6�VoYuvK6I�߿q!��ͦrR��?�����'rKF��!�2F����5N��s���<Z�N^��/�<2�G�.X���P���˙��Vǵ�K��Ϗ�Ќ븄�`Ѡ,i%���f΁� ��,6��R��W&�Ŕ�E�����&'�-*^��*U.�/���G�H��:z:c�����v�F��r��R�M�v�N�����w����Db�� :��su R�ơ�'�K��E��Iu����,�~�P&��-�X�o�<�&h��&�;]+���u�H��<��e|�8Ƴ���$N* �s���j9�~����M��y�{ґ�_�����_.Y�O��O��1�ׁ�M����?�m�y��t<�)tڍ l?�X6�P6۽i��e�#�o�)3!�W��a��V�M�D��)Rq��ڟj\6-�?�V��L}��dϤo(rt.3�������:���ЯM;��p�������9����`Wd��at�X����;&4�-�Lj*;�h�}�;����O�_�6�h|�b��W���`�����Դ4eoS�!jb�"�ɟfs>Up����[�SV��@n���2�8���(�^�o�3g�@a��t��u4D^�Y?�O	Ϗ� ��RzD�~n�f)��W&��ƪ����Ǻ{�Z�DCQY�����GE$#��]���<���d����P��d'�{�����>���}^�筗�=��u��{�s�<س&s�z@�q�`AO�/�:����#����ƾ1l��une璻c��+jv��ݹv��{�ǖ:�I�Tc�"���{��.�k�*G*G*6Fn̸���(f��G����4�1@��I?�kT����uZ	|-0'��9�m|�a��ᢦ�|�#r�#�"C-�D��3�0Y4��`��J����\�g�z<\uw���%����M���W��ܙެ&�p����9�ğ1^+/2��b�]�����&�br���m t>�C /n��a��t����釂��W�sH1��mee�����k������"k�b��&��BL)I�'��k��b��Yhц�o'�b"����\������qhB�J��a@�XBn�j�T�J񄔮u�����/$�޺���(����"�pL�/�Vi�$"obգL&������70�c9o?E�t<��D��{y�-�_2B�+A��4*	�M5!U��U�����jf���/Rc�A1Ld�"X"|��#���~5�c��u"=!�O(����]���}��\T�
��N$q^&��E�%�
#���\̨2��C�1u�NJ�{�n�d�.��^�@����}%�g�^��~&� !�;V�bG�0LѻW�C�KHSj������~ʯ,orA)��0��þ�$���	�B;��N�G�~'��d�aL{�Hq�ڹ,���P�+�j�j.��R���?�;.&���RІ���۷yLg��U(5�*n������3��':��
a�ݸt�3�Ԟd�&�#�b�E>���e����v�B!`�%(�r/���r�3;�nr���c��$!�:p?ӗF~�=>>���U�)�`��I��~������w-����}9pᗡ��:��EMo���'3*N�=A����� ��"�s��&��r��h�'$�Ø1�V�	�ʄJP��ޚ���'(�+o�1P���pc㕦*?�m���X}[����| v�O��&�Ҿ^���^�Y�t\nb-xlw�p�����􍳩=�ō�V������	J��Q����U�<H���,*�`�2���}�>�&<�:/8�Q`��s܂�z%o�N��R�b��ЫD���7�a<���g���#���bf�����|:�����YEL.��(��~��,��fΓ=�.�b���Ƌ�����)	n��M�(�HŠ�ld?5�bl}cl�!שR$���}�Н�^��Nn�[+!��LxZ}_�~�U��U�]'Q�ƣ'�]QϢuP||S����p�)�)(y��(x_�- 3�n9�y;b�s��0������G��*䑆�4��\��y��\�_�xlv߉p̣�bc���ӧ+���y̤#��(���3	�oҫV7�׸�[ösnQ�b���֭�YY�LŠ�1�KX�8~���,����Ezkn���_Z��O�/��3�(���z\C;��ܱ0�sI�#E�	��V�wh�B9��?&��tP0�?�	yL��ɉ&6�Z3�lrV�����W��e$�>�*�sg?������پ脱�#G6��u��e${IV�֐�3��i|��Ȫ�n���;%Lv�h\�=2���{�i~�$����=��T�[q=�J9JW��:,r)�˹���:�&EF	vs���Osw�\�mK~�d�On0T)�<�%���0<6O���c�� f*I���mL{+&������S�LcI?������	jq�nQ�%��#�l���]�d����ܘ�UX�u�}�����;
�O�n�QN[����?7U1�T��D0ڨUp0�Q�P`�S�ۛo2�{,МH;����ų���I�6�Ԅ�X���]k�����I�	$x�|%}�ki�d� &{/Su'P�ѯ�+_-˶�B�����r)ʁ�$9w*��c򟝜h���J��)��-����ZL.7�j��5.6���zJƝ��|��9)��	�D�O�XV��vb����'�YZ�Qn�A3��GOL���^J	?�m��y���ى%�k����B����Ŷ�'�ʛL[�nَ%�Yc\���k�$�N�C��En�oR��'���6���4��F��xWP
���x*�RMY�5Q�w))!ۦ�|��V���*�cOp$�[{go�N@�M{�O�؎�ib��W�Dj9�wG�1b=/qs�;�u(���\�~����GOH�8�t�?��QI�- k}��D��Tl�$�kMM)��W���7�`ҟak�ZR��[	��qf�����4`������X�6����t��~������H����f����j%н�=ֽ�l���}�8Ĳ���O��!���m-���*�����(Xz}L���!��ర�RK0���l�R��_ܪ�Qq�LPW�}n6r*o�+���g`����>�m�`�iI;V��|�>��.��S��66�O����+�^���]��e������p�-�m�	������lł���0���(����$� TE<ҜM�S��c��n��x���%.$��ؕ}l�È#��mD�ƆômO❰
���hZ���jٳ�9&}WD��B����{m�����HF�?l_�_p�'��ݓ��x�����{|d�֋��Qу��n������t?V�Qa� __�@;K�q��[�K8���΢��ע�)���A�j�� ڮ���z;!8*�9�͔��	�t�z��S[>l�ā��tO&��:�j�F�OW����N��Z�u�E�싷
{�Q��� V5���m7Wc��<�n�Q�o$�����������ژ�нIu1*.ȋ0 ���b�S�����B����Ln��<̟�s�C¸�lCG�I�ku�洴����b �p�&����]� �R��H�:o��:�mM��?G���P�:C[6`������\�V0�)��BC]]����W0�`2��p%��b6�L%��
U7尛k�G��X#�݇n5�WP�]�^��Oe��hW1�TQ������ŋ�*���ϻ6p����Og�h�]�jZО�(��{��^��nQ{$�<}�RKӜ��8��-~�Hs%@�" �؀ln~��_�i�NUUn��O#蔖�q�E���\Ksc����������R;��1�\��zaL��yN�\��T:�}�^F���Ke0L��qs}8�xgC�R���x+�Q�>�޼M>X��^���ܖ��Ϲ��bA%�mP�	���R�����kZ��>��r�EtB�%�cS��łI�k隉��}u������s������4.J��!5zj�mjҚ8FXoʯ�?_8{���BI�rd�}�e�눛��֒���5�,� ��~7ġ�p���'B#E�ï�H
%�N)7{sd�t�!~҄�mNcT�d�ׇ���r�⪪�ህ��0���N�������'�m��S���檻0Ҡ� �1�_e��@	���6�~@]�'���`�/�����[v�~OJN6��n���m��������U��Q����K�t�ä��g՞��,��>ϡ�[�ՙ�+�)��u��Zƛ�!�>���

����0�#rl�O'�%6=��k-��ln1D��wߏ�����^�Ȥ�n6GV�0.D���k�g��d�f%�kn6����|�A����;x~��BT����+��f���Y��z�x��k�G�̎�w�n+��ɰ��-Mr�ΐ^�u��VcDA�����/Z�2�A�Ң�_�SGL{엚rz�f�����5ʽ��lOz�^�R������묯����w��yf���;�.�} I>���۳����-,,��Dh�/4�o�#t�7|t�H<�j��O	[��fZ�..��btX�j�d��9G�i�����ӿ=�j�[���)�������W���6�ʷ7H<3RSSWF g[[[%^�w�B(u�H�et3a
����ʛo�x-�`�ky�i��E,��xE�UsyqR��X����.��t��ǭ�x-�nt�fK *6�j� ��CFgg�>q�����_��*���'1��{<���κS��8.��RZx)H� m
��Uf��^��H\�z�|�n^RW5���Cp��A�����,�1^rn�����o=�v\���<��Oe����dCL��U�|��N���c��D�BA�����Y�[��A�V�Bڷ����������_�Hf�ɜ��M�b�BHn��oq������9��`Ŝ���QF��y2��3=�~�3��z�,��$�s��w���I]�l��22<,_�X�˥ߨ�Ǩp�z2���VKCg�����.¡|��s���c��y�I,�8:F����u�(iX���2�2=���CH3�M� k
߈��kj��EU9R`��='y�����P��e���Q������S��C"�÷pm��"��)��^�E��XÈL����xY{&�z(��/�@�r�ѢH���C׽GQ燙���yi瀋�֬Aq��9��e���<�}@�i}�>�[�ī��� ������de�MjK3�N ���P�7��P���`��U��x���N�_�UD��jj����������Ϝ/��	7j�G^���.�2,b�2�d�kPlJolL���mL�����ws>v
b0gz~I#K@�ҋ-j���nQ/<=�[f]��t��)e#tF��r�|9�1i7_�Y\�=0�aDm�p�Ս��M�NT�k�E+��-�x���t�{�/}���������B��':�,i�LqQ��G�H���h�2��� �;H�8L�J��
8���{Lb�������}�\ٝݍ-'~r���z��◚�X/��1o���F�ψ{}^�磍�����!�I����cű
&��?=A-�7��X��x!����)���Y�ېfA���D푙?i�;����;!��Jm�
9�jҊv{�lA��bjtp߂�xC9��kW�lG���K}�d�H��Ԃ� �9��ѣ���	�܇e�,�t����F'K-��22�ҟ]W����>��0ʕ�)�M���B_>�B���lÈ��������%���e�a����N�.��:���𝞼�W�|�[��xRfY�e��_�b �s�z���|�D�gk�	���Ap��]���Bu�����|חEC`K�Ս͌Z�����;�jq�hq�z$�*�4fZ�G�2�2ii�Ŋ����#/�\&͝58/^<���|y/_�W���m8�eG8u������,��kY�2:�(My���4��v�$͸{�������-`�T�u�/�\юl� �}@�az	��������xr.+�ȡo[2U����}R���A��!D&�!z^�Oܛʓ�ʊ���q�̐Ʃ���'����7�wVc�5�y\�m|��V�Q�i e��/Pj��x������t���C7ϡ%�O�;����Q��!�kb��a��+���mo�F�7\~JF� �U�=I�_���/�&���A�����`��?\6޼O�o���u�ten�Ҏ �+����]��`���.Z|�/b]{���э�]�K�~��i�_��o��51��*��>�6�O��q&��L��>T �a����HP�sB�������]v�s�ϟÚS�'-�;�'U�:F�I*�����~������z�B\����J�ka[����!�[��D-�Ȅ }�l����{r\�7[u���Ð�!�q)Nx�|*'9Q�8n#���%$�_k�#�5�~�"(FE�\n:�(}s�s�!3t�1^뽘�)J�ii��Z��9Q��*FX(:��,��x��2�	22�򊯺\f��_Q��0Y�P�2|���-<��R6�S 2b��֊�|U��V�2��2��%�*p�Ĳ�afǢ��� ���CCC���5��Q~�)%�u��tL^��<���x�`6 %�k+�-�,-͕�jLx�x<%O{�w?��G�$��7�����T�R�ٛ�t�Q5�,S�uKV��i��bJ��Q�6E ����� ��m���B'Pn��)��3H���@@�>|��׶Y�.���^����گ�{MkX�=�{�w,ɛ��	�ex|�zy6�DA3٧m4�R0��F���FohJ�Jjƶ���ӟ!��������ߗ|����0��->+hH����)��8�k�KY+��0J�d��3>���O�t%��j?C�"�7m?}�򌁟_�\�րә7�Vj��������T�k��>x~7���Nx��0R��.���Ӊ��ۅJ��/} wtToK<`?�a���Ą״�m:����yMW�Ź� ���������9#~����ڴ7R��c)�����\�垐5�Q���Y��LNJ��ح$;�/�>Ik�� c	���F2��������C��l�lٹ��~-�G�Vx�Ix{M�^��s\�_��r�U���66|�Ϋ������}�:����dLC�igZn	)�N�2�s�������)��4��e0�d���6;�k�_����0����!��k�F���1��k���H�����R�N��f�


�����K�[K����
�s��˟�
`��<��m
�a^�j�PҠ3��~�t��ŋ�*��� h�Z�����Ͳ�z�AB�CP�� �=�т%+S����-3xN���l~�X6\ ���x�Y���6�I0�La�7��Db�;�k�W�zVYlw*����33�رU��H0t)-��s��|���2�Tx����詐� ���7�r��Ӿ��Y�1���~�eo˰���!���|�d-�څ4Y蝑��/�JÉ��\VV��xS�m���4�D�~�Dm��>��n�#3_8k�C�."X ��A��erq�ˬ�e�׉$�KN���۸o�1UY:[���5��~M��;O�������M�ƻ���=j7�

��{0�o�~!�-,I��"G*ʇ�/_��:�`"�kA��CJ�!d��?�15�i��@yTw~NJJ╫:-C7���~Bk&�Ğ����4�g�(�d�OOg��ED��V���4�Ʌ�)_�`� Θ�dm�m���GǙW���T�����2�MH�H������9����7G�7p�%���B������ƛH�0�eZ����*>���[nl>'�`�=0��39"����StE�Ϭۢ�SC��&�V�;��+:K��^��sb���mug���,-HK�k_T6�jA^n.{o�R~ ���khی}n�B�˴���,�"}�>�f ������>/��N0���R�cM�����c��n���qcY�яQ�G������4����]|�>i5�^�;Ӏ�z��q8���&�:�i<1� �㼸�?ߵIƋ�Ĕ�g	�)^8n�l���^-�Y��Y��#O7�I3��{أ��ivc}�x�b�<�5H���e�2d��+3�>�2�i<�@]��Xx*�_��ml�	9��m�-�$9�� _�׽5�����i��[L�MM�7�
�,��'�8��򉗻�J`qkE(4����d�Ӄ���v�w��S�=�6c�/��5�m��b��2;<�Fj�J|0]v��V�~�w���Z4�6d�T:�E.^ϼ��]F-����3ގB�u�q��V���#��駪q�HI+~�~�R���а�k�~p�~����qO�!ćЇ/�=��&.��̓9Ξu���#Z XS�аF����Z2z�9T��[[_�T�۽ F�2����3�OyR���ػ�zYd[o�9@����%o���r��z��oj�:?
�O��3���A�k����y��K��^c��q�3ޔfff���u&�����ze���/��8����F�0�wIIb)-k[m�s��S��s�]��\x=��?y�!�̵���D��2����?{M~��΁Q��2�<�ldhh���|�P:�aK�kF�Ǔ"4>���)�;��Jp��kM\��B�U8n�:|)эibjs��dz8��jG�qAw�M-Z���a|t��6�s���i��|�������2{b�Y>ټ�n����fJs�l<es,%�~�)���q���=܆_ѝW�)��;���x�������
��{�����ɺ�󩏭Oݣ��+;�՞�ͥ�ر[��;D�ƫ��o3G(�	�T�AAA&FƬь��KBڻJ�PÑĴ��QF둲��tQ���K%���T#q5w�Y�f��L���`֜���$հ��&�����k)�S�˵w�5��)���D����Z��U'���4��y�����19%���$�<☼�˚yzo&�yϐ���o���P�~�}��r|�����"�6P�]�*#{%�ޢ�Y��)=���#.�������=+^�l�2��Y����U�9J�Ϙu�A(�h`��:�1� Ռ�u��X>|�6�cF��_}�%w�����,h�� �g��oSS9������%��!ܑ!�r��KI^M7��������)�i�H�5��Y7:nv<~(ZL���¾}����[Zp7��D_�=nue�9���ɀ4>��c:p>W#k�Zm�,(5��3��.ԙ}fE���P�[���ʁu�^:ʒtGv
#R2�����6<6w�l��@��;l���Dl�L�eF��G3U�HO�8��Z	�Y�}���ų�	��8=���K[ߠ�k2�&�s�jVϵ���m���E��˗�����u�R��N��C]'�,��CQU��%S	��a;�� �W`:^��L:ka��+��s�!!-�h~��Ӛ�'|�L�5��l48l�?�Q�U��j��yuę�&�>�Ȣ:lN�YV!R����7~u������n#���{��xg�����Օ$Ag�|����Rfo$��AKr��7�qR�lmm����@=��-�`m���?��#Og?q-���d2ߨԖ�p{bu<͈yyd��������mJ�������׺lzi<@I����B��SS���BK�K���Di}9���VH�������	�W��؃�Q��`�%sai�����=xܳ+v�T�
�L��b��ل簐��E���|���,��X���@��j�N%�4����t���sթ�;�'�n汯UԨP)1���h-��}<���{]N���qn������2����K���~-�����f���egV�W��$Y=Җ�������\��� �(�����Dt�ي�=����Ys�!�	�����,��Ũ S,Nu�6�h�>�B���)-y|���{e�FG_��JF���G'i�Ěy��ԌU�����k��3Yu_�J{�;C�&�t��C�';pPF��B������h�i�ō��y~m��#��=���ڑ3�$�W�وP#σd��|�e��Cՙ��Kk���t��]NO��d���d8���p=�J�$�ϵne�}��]m��6jN���}��l~MY�=�Q���P���˼���E}aǓ2!:��O�s��ͻ��ʠj�@&�+�~(����9��Kd�
Y�$�F�Q69QBJ�'=B>���q2ac�Y��)s��}|��!��>'��O��"L�ê��[�c�G�m���S���3��Ůk,���T&�4� �gÄQWxz}��l6�׼�����h�^(d��(�h���W�l��裻2;$#��g�@
��c	���N����9�*�l�� ��)�{�:���p�O�I#�t�����,,C���<@�����g�W\��A�)?�|I�2op���k k���Բ|�T�M��|Mx��"}�=̈(�2�aW�x�������+��8�o��s�!N�5�|��(.�����5����n���m�Xc�\�pHOK�f=�s��cNn���{�u		��J�n�-,MuA���|#q��'I�c�(#�K�/���z&���ߪ/2GԎ����Ĉ�n��I���J�vG]?�d.!H8�c�lhoo�����I'�� �^�#��1���i/��m`�kYj��	��p�&yg!!��Xb�~��}2��{_ǡ+�{�r���p��W�n���FP-?jF���Ĝ� �]~ɨ�;̓u	]{ak�B�߱},�z�>��������edn�`&"������ U�EG�qb�_
�9GJ�#��s=e�F��ÊN�j�W4����б�5�#Vr" �7#0Q�k����w���l����цh���cc��lO[Ϛ,�5�z947Ɣ����V�K����0��ʳ��"*o����ܠC���/��[���
�1;��=�i"�u|rCs�1<<L{9����HC}�0��E�Tv?.�$�?Oy�o3�+n�[����ț�i{�m2 n��Y7����p�㛜 �z~#��3gc�)��餤��9&�z��t�:ZR�V����G�3�]��;:SN�R`��^t��������s�	�Y]�)-�nnnD�C!��:�113S`�5:|OWUU�;ƞ���)�0�I&Ӵ��"�~�g��d�bPm4�0|<.�]c�C�CS}=ǘЇ�w��ȓ!�3�[9a+��ؓ/X|����=���6���$������s��M--#�x'QCta7��O�K���ΑkS��ODD.^�(S���2��8�НoH���*}�>�3�X4�	��kϠ<��J��h���+�<�Y�[o�d��'A�Ae^���8住��mt������n����)r ��D36��CXJ�%�ȹ���M(L�`: �OJ���~�?{m�gOc#��//,.�g<R�L���Z�^��j���'�cA��m������Ջ��P___��56(�(vW�xNU��١�͖�sS���F(�.wO�'�B����7����3�<�4$,3����OЍ���i���� �����fV�r�f�9�5%���2�A��T�&Y-�e�h�ވ�r?wb���F;b
�޿Ő���BMt���=�qYY�х�i�*@ƥ�N��Qn~��큨P��Z��ˢ���qRҘI
��G�_ �##�c���7���W`���4��W�$�x��#���f|n��˪�J8]��h���J�v�(C|^�ڶ��jг�y�����B�d��v��
G�N�T��}��ζ[I5Rz�]z/�n����
 �s�c����}4�������d��g��-�A���������rv��U�;
Տ��A��9�����[Ǻ��}�k�%�����x�5v��7�ᚐ��A�����+&����L�<JByͣ�@����C��	j��眢�0�#~l���#�z ����)�����n1q[��H��E���u|r��c��Vp����G"�+q׷�k��:(��A6,Tkn�ύ�Z�mx�����ш4�H'rHt�����9�@��f2֞_��t`��nw�ˁ)� )�LL���mo׈HH�������N�k��?Yq4�۸������(B|�n)O�iJ�vqBE�>̽Ш [9p��4xA��r�횕 �C�&��O`�����N�5��H1�w] ]ݝg�Atf򵏵��b�x-r�c��vŽ�N ɁG�`�; 
$yDhހ9�)	���7�|:h�����r���k�=E�]�QR
Z ��S�o���Y7���Fq�ģ厓��X��*���Z�is�;;���@lR
X�\[��﯊H�I�y%}d>�Ň��{�sOr������3COOLJ°���T��`<�+譣\w�q>EO��L^���G�g��㣢���3��!D3��&�l�/N�q3��=��*�6�47����?��{�Y�Q�ڔ����|PÇqt��N��@�5uu�wl��d>}Y>P�v�9CV	�D~�y8��̰~��8���/�99�	e��t}��w�#�D/q!1h~���3Bo��$�P�Hlll��M��}� 2P�1����m�(�gGF]ݾ#~ثAV�u��Vrŏ?�||�v �%��oT�Gm���߮:tHoq��p��8��b�����uu}�4��YH���u�d�+j�>;k��`*3N�Ԗ���uX.�3�\&*1�#�x����x:�n�������|���9cV	�1vB=�J�8TL�b ���3�A�@�ڽ���-�WA�� Y���wo�J��˨]���_�l�TR�]�h�			�D��my�s��$*�X�rНp��L�3V:-�l��2(��_��*���q���رN�x��P#DD��\	�>]�~�A�����-�lH2���+@ѝ�w陵�[��oe+����7FV��|�1ð����]x8�9�A�%����x�}��0�iq������0����9�P�����ysG�t�ɓ]5z�V�}��QL��
`�g�/j����Ȕu!��y���I)Ǐ�C}�XX�V�Ft�|�ʩ��C�Cz���"L}.���f/�������3V���թ�W#�m������J��b�s�D1�m(	��K�R�� �	��3�,�q�cc���F��hkBy�?��� �ş�y\f������w�sǓs�?FlHA՞	�z7N5B��N�R�C�$�rJ?b� ު=)�nrz�Z':c�Z�gW����J�\�.--=)��[9��J/w��w���(��#�X�i�_~GP�+!����X].�����Ж�'{ж���5��-�Kk���[�kZL�p�:�N}&ˎ�ˮO:��+�<�EFJZ���Q����S�*�	�.�%RT_�*�I�}��!w�ڣ�E�lu1�0I��4��c�DC�JX�Hu �2�SˠR]h7HA�����ͻ���|��c��O޺��q��-%qb��O��JG��҉E�ռ��X�����k8���^�#{+&�Į�� ����J� -�ڮ�̟?s�C1�5@��������y��
�K�Haa�z�J��k��:�{�٢��^(5
Vx�����fӄg�����)�c	1�>1Z�Oع��@��М��\BWƂN�:�ݑ����t�ܹ:�gJ����9 ¿�������r�(�u�s�=���Fe5:.Q=2�KI@����R˫�|XC{GGC��旕��tGWz(�u�<��(<��b`�'0���RP��sG���C6X��g��S��H��9�_���NH��N����L�WP���q����OM�Ał1�P��!]�9]V�2�+�u5�G"�\T���(J�U���妉KbVl/��h�v�Kv	?i��/"Ym�*�]%��N
��!�0*��L�lD�UbT<�������'�QS"�����-6rs������WD�Ń�cM	�_ �PbO��0#C���^O�b�6��ţ��^�xFO�3����N-�Qn=�in��$*z����ĉ���/3h+!X�|=�$�sdW��8�/���_��D����z-��P���Ꚙ�f�����@0��4=��'7����~��Hj�F��R�A�������ht�V�(E��X|�G����m4ᮭ��3񮯗�n� ~1t�U4�koL�#�mV�6\pvmJ�?S�~��eٓ��Q@A�U_�F��A��_�d#)�Z��k��p��=�4�1 �9|���F������+xy�̶`34��zD�&_�~�]ܯ��|%t��NJ8?�C�|�E%F�v�-0 ��S=�4!�AA�V��C���l���abFX��\�^yCT�u�ۻu ���c!~��������|��mj�|�C�m��-��=˴��d}��֎<+��0D��]Kj���2�B9-����G�D1Y-�����իW��|Gِ�P������Ru|�z�H:�rZ(V��nQ�¨�� �¥��yVr@PZ�-�c�Kݏj�O�_,�q|�G�Ca���r�/��@I*���]��6+��F���L�5B|�K�[����5���Ͱ�y��4��j�`���W3�ޯF��y���y�/num��)<���ϯ~���	wu�򁭔����Dd`+@�o�.܀���`I[�޲�5R+��Ԧ9�*gm��P�����X�>��Q��W�T�%��A�9*�v�A���Qů_e��y(�+a3��X/����?�r�I��*I�����0���;��e��+������K�%y�n�w�ܓ�=��S��wLLL��6�+%7B���jv�4�4_�1v���2�Iq�C�(�ت՞e��h�SN((�(����:nN�I��0�0i�
Hj�G�Z��h������Fm�pJ``���Sg;2�����7_ؾߑ�2�ٖ7B�#sz[��`���'����(�ee��ra�º��� ���G���-)ö��-�Jc�~ �ՅǤ��k �[��sef�2+��6s�<ljj�v�N�1�c�[~�M����dy�%+�`���/	��4��z�iM�V,��q��ͮ��~��U>O�5C��V�m|���|����=�?��19�s�ZrTRP��Sޜ���N�6��T�z=e�x��F���|�/
�(	����~R�Ь�g���:<��F��wxTwJS�����ש���$�n+�(~���ӍP?�c��&�Bi�����-��#�	����<Ǡ�趝Fr(b7@S�s��T�N���QV��J�6�&�(���d3�b����d���\}�S(R����9ȜR�O	�5�[ݘvLinV�qœԲ�Qw5�C�լ��(|���& �M�9 1`�������ث@%�v���؇7��7�g���.��;�U���cĜ%pC�]�'ʽ�b'644�ՍZb@�����4�g4�#ٙ�W�t�>A���^����w�%�?�Z�շnbK�N����HK�dy�Z��������Eս��cAq�
�}K�;+vB.Ǻ��������!렞�Ki	)�UA��²ZB��FVhE4N���@�9�ҟ��\ʲ�F�qQ�STT(���S���t�+W	ԯL����.%|0������ORQ5����#u%u/��+ U``22�����_�����xG�rJ-I�#�g����������8B�Io��@���.�����EGІ�����8hN�z������N�<�]��� /�k�(�#o�~)_���#q4Y�k��#J{|C ��m��K����h�
=��z��� @ę���ܺ��z�GbV�m͕*%d�i����|{{�|�����h)l���'T��m�lB蕇
;j�������]��)�ո߉C�x���ʞ��6�H�h�:��f�4��v�և.T��ӓr��7__6E�٦@b�T�ʣ�mŗz			C����$��h7Oܛ
"��a��Q��+t�b�;_5��˖q`R�����˰R��u�����d�\���s|������\����������O��Dh|ʴ+d���Q�OJ����+��29è+���q�?��9�L�`yf`lr��q��%=r?za���F�����f@@ P�C�g�N�M)�K�����/E�x�k`F��䌇��,��4 bk�p��ݛ�S��#*�v|	��b�����j�ƛ�T>�{N�D=�d�7���ߤvX�V�r"Uy�	Z�ǜ�$'�����ӥ3��J����c�XI���k6ڠ!$��z��Ot*�>;.���`��3�̄�@�C:����@�t)Z�^���
���'���!��q�U"E,�I��� Hх-��|�v��]4����\_�����|'vj���6s�פ'�R�-_RR���4�����`>�~�?�4�]�v���x`��."/	��	��� @��"R>�� ����F�Q_�f�FuЅ��qڿ�Y�#����w�F -���&�9II���鹌�����$��xy��̊�̀'��]�?Sz�L֧���LV���ɳ�Om���Lsr-AI�N��Q>P(�e؞~-�KL��)��T��pA�)�4X`��[R�@
A	��–��OQG'6!1Q�0ܤ쎝�_҇���JJJ�z=hioOpvv6��"wNHH �w+�l��@C�C:�Nww����RHq9�,�q_c]�^ZK����0��q6����4�O�Z֛��Km���B���G�'ڜ� ����/w��5��$&$�fs��:�2�UH��'�n�B5S����QuM͈m�C��"l*�n����M�ލx��ɢW�WI���<����Wkn��;8��u�ڃ=;>�:}�@ثءm�H��ڔ����sz��r%�@�R� �B���C�bo�U�d����K��N&%|~KNu�L �:l��<����c�_f��䱛�;̔�RPW�W�V7�>�_H�M�^Bv�2�s(�PO���܏SN*�,�ߋXv[���T�?�g�_A�y78NEE��۷7  .^���Õ��N��;�N��.l�:�1Z,�aʃYIPŀ6��5���B~oSR.HW�?011�D鞦�Ǥ	pi'�+������gY_"�5�Rd���䃨����Ea���G|*eRB��X���B�(�Z�M��`�_G���D��=x��L��	9��6P���^%ˤo�᳄-/�!r��Tt�� 64Y-;
ʱ��06m�A���}�e	v��1i5��ߢ������`�b�'b�;�c�9 x(�����t���!�<� 8�v�ѡ0D� ��Ы��$"�k�_2���>;T=����w'�*�i��1y��l�ϡ�������74��#c���J�;���:0֔8 �5�9e8DO���'��ْ�a�\:t���7�C�|��R�/�@e$�<q�壘��}UZ]V����"WL_�]P���..g��
5uttZ�~Z���Flfs�7��E^E��2���/Cf�OK�/-��~��;Z��q�5d��;j9EE�����~���_%���A%
L�d*!k\��U�{J>VS�J���jEb>v��3���j��0EԎ܌�����pVf
��*���Y��ݩ�<�߾}[ Q�*2N�*�Y���uy�k�5@� a�J� �H���&/[8�����/[O����aWQ.(Z��Q�?�Y�%��h[�r���oz��h��'#���"$�����UODzmģ������,m���B�/��|�D��|��Ѝ�b��/7s�ߧ
~)o��H�t�{��@XĜ���T����4�໨(ZTa�|ka�bi���zrϞ=��FA�2����L��L��4�F��1�r,ʯ2�������>��蜝��Mpp��Q\D�'�Y��k�8�M�Aك`�0>��F�egy�=�0A[EWQ�C���Wa��~��c|a�˲'��CO"P��������{��	���(O�C�y���߉���=������P9���M�T?RRA b�3�YA�>BC����T}���0�4gi��LEz�J�|"��LWW��S��UEw��*�o�9�'e޺}�'R������c�B=yx�Sߏg^��
`�s2C�jc�h3�L�+b���Z�L��Κ�!�	��T����������B__������:R��"+�ݷ�1��y:��31� �@l�HM��������w���?7y����4��Nԕ���,�n/�J.))�)ݠ���NI)aӫ���x��v�5���]�e�3�SU,���}h{�����z�y�������1�A�A���} ���WVVFg��1j���X��`?��u$a���:�ہ7cIv�3M.�6H�x��'0�Q|�yF��U�4D�E���`	����i�����<�Gю;����V���(��9�`�P.�����ee��b�-�ey�c�A���8�3
\:66��`�5�G�X��|l���Z�+� Ғ7�iF����������I(�A�>�rNj�@(����u��R�$�]haQ8�k�-~*�0@%�V��vL��h	x�X~���KJ������8^�����Bj�=�[��~k�����^�Co��"_]�@t6����4���՗��)�W�K5���fc�`f�h�Л�ٵ�LR�4�ڛ����3C�w�x�@ر�x�X�L;rV��+� zM�T��'w��˗��9���t�jI9�]z��X#j�(�O��������=L;~r�]�Ә�e��)%��v=�Rx8U�#㸞=��d�@� Rb���^w���%�͏��g3;�p�#c.�-%��(l�Þ<م��+���-��p��O�K�S��$��Đ�Gl���ag'�u �����\O�^D?~�3���C�^��y�������춝��	{�'A��qff�׊���&�ik䋼)qV6��M�������.���`逷�"��\ꄯ��羧!��K3��e g��O{�cW���߬� ua�ʁ�PiA�����v����7X����*:�B��J��yYL3���3��u%Cm���ϥ��W��������:ᗢ~C[�Dr�Ŕ	���iء��,��a�V��z��u���P�s�)�,�P���"�8�.��Ѱlm�0E��c{-����y�g���N�$&��OOK�^{����ma-%�|�ܾ�{��P�M%�`%�2=''��R��E��'���
���F5�Qt�D`���[*r(}G�5�9�%板���,9Q��������P����HQw�4��X��iӢ촐�)�Hd�6��:���D�۠���"[�d�B���`"&M�n���}�������������s]���y�s�s�攚�e �'Nq]�ͳOJJ,�`0V��8�&M��S��wϟyׅA�B���{�H4��}:t2q�5�uu����7﹤�s{��Ś]e�{��~��܋������.�^C�O�ޅ�}���C��?��ߋ�'f��+ݜ�?��
h_�\|��|���,,j�[<�t��F�o��׿���O�P�I�	���
^��OwA�t����"�|V��{xb��i��N��
.�9��]�>~|�}L��-�!g�B�|	����q�����Skk��}�i�������;oL�>D��fU�c���p���"_±g��f��K ֑����޼A���B�I7��ߵy�1���M+�x���s}vh�2��]'!q�̻�|�}JJ�ϟ�rL�o�_
��=��s#Ӳ$��>��$�Dz��mI��p���m�>�:pP��?���.[������~����As�i��+T�Y#`�Ho#�j���/��W�������kfM�Bs4š:7$a�����#ϓΟ���7�Zh�e��?��4Ȩ��>ɱU�
%W�pGY?wh=��WY1̞ff�V\=p:n�=ڱ�н����Id�y��|�zB�L{��$�[/2�t�t��+t�<k��u��eK����A N7{ʰ�) ��`�̥�{+%))��ҩ]]���/aKu��~p���W�*WC��(*)1��={�2-��q��2?��{�n�)�$y�bR��6�h|_�숊>�A,+�mdl�g�Rǩ�b���@��'O>��B���3#�%�����R�"dn���mϐZ$�<L�T���7)�j��><�+�ܵ�ӻH��?ʴ��j��z�/����4$D�	���v�+5ㆇ�;���_U^��ڟ]�A&_��
��gӿC��3����rh
,��>Ϸo�f2�6*NxoLE��Fv�@�8S��,6�[��NU�d�+*5�T�6��Ǿ���쮧�ѩS�������o><��)t/����B�f��-cx��e]OoI9��9��Xwp~��	_M�I�n�);,�<�����3��NΛ(pd���i#�(U5����l/u�cf�)�Axe��Nq�[Y�	���#k(�V�v��\V��ٴ�Pߡi�aYl�b��;3�ЪȕKh��u3�\M��E���χةCZ�_�~���ϒ�`i��/ڢ�t�!eI�?P&���%��̓dOC��n��O�d�]�Ç��� ��T�sI롛7o�}?jQ�~4�<�[�y�҉�CO�6�z�z���Q��FC�����>��=�~�a�;���^g��]�S�~vV�Bt��|�QĆӑ;7[��9�b7�����1�Q�#�I�9g��]��5��ĉ�p����7G�bb�_�Pܱٽ5�3��rc:;{W7c~ݶpv΂B�^ZZ�"��k�Ii�%T?;5�R೑��"�FU���z&;�����bˬb�Yo��>>E69�Vo7���M]BB�_�屚~���y�l(�� sG������%��]���}������\�Bh����EP��rAn�~����""��3-B*m����@dN�U�g��q���P�\h�oim���˽&���T�.�ϖ�H���[�O�Q�ir�h������p�����:��A���R��` 2PRp��682�ao��~����<�ݏ{�5�䷛4��A/�;*�Y���,_��6�/�,dMZt�O�c:����ʭ

L�K�i�:�'���,b����&�S�E>EE�i�Qs�_�L5`�״>2���l���_{��;�TAT��l:u��w���@�uu����N��P����_8|�S�����2�x&���
ܦF�F��]ȍ���H��]_�7�Ե���,R F|懶b��{��rЇ!{��~Gh󈩮����C��_mf���W��|F�<c�~]s����h�p?�W���O��N�������eq���b��5��zǻ��(6����%�$^Y��е�W�F̍Wm^�����q"�H ht���F��X�����U:hB{g<��|{i�z��fDZ�Hy��f��l�r���,���F\O��0vY��/�S3(o�\��\&y�.�Vj��Ϸ��ii���L����/��c��Ɩ��VDPh��
C�Y�l+P��I����ݲf�(��{�U;�<fD����ŴިrZQf�s+t���^=�l�*պ�T|�DMU��Z�,˰n׵�þ}Pୠ��n_=�d�\	}bD�e����I�[x�p�z4[-#--�0S�ٽ�5����3VV�oֻ��m,��,+K�����Wf�9�����g{�f��x� MK���5UUC��^~F�Ӄ�� �4{T��8�� {j���.���_�=���Вl
}u�e�ʯ�,4ڱ�MKK�6��v�J(�˄���p�no�b]ج6����:h55�YU.t��7*kMo��j�x���ܡ(�Lh��jv�N�b�����}zb5�C��>."x]�͒�\�&kkk���y�ed���S0�,g�%�r'ؖ�,��N�N fF���>"~uX�5�kѽf+��Bn�,��5������Jq�,�jr5E:)ŮP9'?���PLD_�Sl�-��J𝬌����nK�,>��ْg?�|��e�������عxv�9�b�%�J�b�@�����0Z�QɅt)-O)�FZ~A�q��MI�������ʗn�]k$����H��;vUGmDS��T��Yi[��"��]�ot�1���Q���*�r�q��Z��\�M=$�g�t[ǌE�agl�����b��������kb�f��+bD�˽���f�ie�EE>+ŇA�Q,U��%[B�|�z��@�������d�-ǾK�p6�[���T��9�|2�on|E�g2)�8�R_���u���!_�[Wӽ�fʍ���WS+$f5���ʻ{� [��	��5��J��+�/;X��~��xz�}�kj*�f�N�H:�;�:�	Z�\�<��=3���/xU�d>�8\O�,�B>э|���0y��jϚe��1���*��N�)0�I t�|%,}��&#s!���T�GQ/�Q����;���\��\,B��ٯ�d8�m6����3�����
~$�W�i���O"	2�c}�g˂��G�$��q����X4�-�l�<�%��|���EƖ�k� 8���_�~��RN����C>m<�B��o����Lb��*9ш�ٝT��	�q�Q���J��ጮ��ж��dߥL%�� ~ii	����\.�=;���?x�(�{�2�������l�x'�`1�Fŗ�f��ƤYE���m����h�tS�K!�tg���#�:��^�,n�����D��v���P�A�
��K=,h�ۀǭ+p�Ӑ�aI��*u�~�q#�G�N�퓏J���jEW;^�M�Hr�K��s{n�J�dv<�R�,:~����s��z��I5���t�.��~��r�
�x0OOŔ�ҋ�L�V�'���dY؟��R�/��������1e���W ?�Ft~5^�����v��Xx3�6�5V 50%��(Χ�꓇$���F5�'��c���%�@�\��G�bl���[�4��8n�9`��jP�El-���p} J����j.�}�����lΪ��S�!�E^2�\Mq�Ʋ0�7+mС����X�%PʺDhU].���ͭ.�gǜ9���-����557w!sg$h����yЕ�뾮9�*fb��.V�&��Kw�6[i���%���Kmħ�B%�vf�3)I�]���~�7��/��+�*/Gr����es���y!��?��;�J�d�y���>ȇ7a��V�BB��+/����S�V�#�}|�fg�9��TYI;i h�D���>,���?n�.yQP ���~aC��_����&�=R��|��*Ò����]J��Gd���L�Vȣ?��.=��}���6��b��w����n���g��تTFC����ujB"K/�i�����G����P{ׯ_?8�hP��^]�^s�Y��?�oH���5�-X�WүX4�h�#���J4�E{����|tl�U5�͐宋Xh��=D��s�F�^rL��l�3 ��PW�+���׋Iayyy�H.�t�X:>P.�Քa6ؠ+�᥼F4L�,�$Z4�Z#�������[�+>{����]�����1j#_XE�)t���G{�#���^���h�2�����^�\
+r�5��?�#:�#4C �h����\yb5�)�zlտ8Ut�T���%��d7Yn4�4�mq��0�볱T	7o��g������3���"��B>�
��j�g�}`;�p'��H�w�����ć��}�QQO� �S�q�p��vW�@˓C��������U>�`^�P�V�!�1�"�*K$ދXB���A|�v�`���^���]Ǭ&q�J��s�����ٹ�����Om9
�.��<�@���=��h ���jAo�[�ԋ����W����ע��T��Ϙ�o�OGhXX�������,'7Wᠹ����\`��3/�1I췟^PRR"��p� �*�F;0vq�7�GD��fc��n�L�`Y����Q� `
�T��>��A#����xQ��DXU�� 
����͍�q@���@p=8��%뢲ɝ��MsS���b9�-AJ"]?kd#>�"����ѝ�j�Z��?ӳހ��YKۅa:`��г"��{����Jk�f�f��q���R���nk��6y,�~��c�xj#Mt`�f�ޏ1<*d���K��C��g�I�h��<�t�P�������U$��ua��0��Te����:��_�ܒ ��ljߜٝX��>V��Z�(Z�X�y�����_�����~vQ�˗������L�JOL��Ҡ�qFd@�C�݆��|�6/o�h�����Mv��l��1�p�
�1�I��6Z�VD�B̵�םxX����DT�f|��I#��r�@�^��y�3r+yK��XA���Nsb&S�2��4,�]A�1B�'�Cۡ�ܮ�213Cڤ�wڋE�pV��ݬ��E���-5�o���9o�9Ya��*��TV�Żv���B���$�pz_��4÷[�+��f���8ͭ�2=�t�����y��g�M���Mn88��.Ls�
�����eB��k����&-���>����,�Zjg��9��!���,��C�`���i����{A���\5%�[�TF`1�CuXk?�/ x]���J���U�9d��f���]=���Í��a���"��-!28��`g�#�0����&g���W��NߛϷ�"�e��&�J���ţMfHJg�N^F>�>b������/���N�!%���uˤ�����[�s�w�::�`���D (!=��v��:&OC��X#�g �E��}}�(�o�'l}D4�j�RW���C�M!��jܐ*��35/��zB�[�T6Q�&����F	T<3����q�=�L��*{�2z!k`�989	ZrB��Sj�c��M��U�[w�M~q�����:��+{R� �Z)c톱�A B�X��Ǥξ��p����xvH��G.��������:}��ę�2��*d�֗�ȤN����W�a�aF}U3pj��_82�Z���-!03��0�e��J�f�;ھ4�I��J&Rg�.N�|�~SI>�	����c���s��A�7�{���ПiQ�Y��0N���|Z1p4�����^�fBZ��6��hbzbx�z[V��܋ə�V�?cR7"���/�rB�taf�ƭUFFF����+C������w58��a!�_��/��N����RȖ�. ӻ���|����A �Ρ����&R�nZ��[�!\�	�eMDx��C������H��E�E1������g�0$�8a�W	��/�]��:�C��k���3NE����xa�Կ�|{W�R�m�߽2,+���(���Č��0:������j��eB�X!� -(_�!��v낏}[����aA:�z.���WW�Rg�R;�H|��ya�o��U���+r�V`o�a��MC���^��V�
YD�b[�ཙ�AY�X�di`Z�͞��������{ȣh���w B�r@�Fŵ1\�O���� G�K$��K|��?��t��X�h����	u(�`�!�Pc�w)Y���s�D�	2���$5��a%>J�VeRHW���G!H�YQo{L�B�R.�g����Ճ���7ЖO��KCw��-�ҡ(��OS��@ 1.ž�R�1&!��)o,�Τ6R��<iYV{	��m�1�@}�H����{��v���T^��:�P�����U�[���@k�Zc��V��<&�_����$7l��p�gU:��a�*�Z��PA���_�DLf��Zo~����{�0� mq5�*[ qM�Kwu��,�������[c��$D�󽁢ET�2-��0&5��}�E�%�l�	�P��b���،��z��h���ҳ϶�C��YM���#B���~uXmd�=�%P�I1,X��|��Xy�"�7�2����BVA#7�i���ۅ�n���?2�
�&6�6I��T���R��s[�?�
���T���Ŵow���J�����Y8v��p!�֗�{:�Y~&��5�6��06�V��}�-��+�I���Q�������s��;N\zCsy��d���߭=�oρ�����!�ϙ���QV'���6{&��c���㥁 ��݉��"U��\j����ˣ�!&n�`��oe�@˽?N�a�I�/QD'�@A�s/�Eh0O��{8,�t�������T
����j/4xX�i0�=�)��;��mr>LZ@xK�ݡ�`5ǃ�B��<U� g�󓰻�84� W�B֝���s�%O��s��w"��{��r���!���>�i{y��V�!��W�F��a�L>�>MK&^؈n���zM��~T�ݣ� �Zh�a�9��=�T�]$<#��\�{�RJE�����!��P>����U�9��$.�F����c�md�Tll=�AQ���zx1�a*��'�>�<#U�<�����r��{�zH�J��>B�~�p�/�"���r���������@��w�W��pؗ���o}Rԃ}�6���8��IdxσyZ��|�����_�kYs}O��Q߁�ۭ���)�~3��H�/XB�v�.V���{>{o#��#%z�סd�`������6����?3��BJJ4\��O줔#�X�I�=�@	�6A���Y(�����7��ӚJZR%�)iis��^�!����S�*PwU6���x>�})V����|1��rix�9���z��(J����-�0W��b!c�R��J3<����3 psMo�#4�t �۞d��m�Sf!��XAyP�����<G=�B|!���E��_Le�6�=Fhm��������e��E����=��{y��c��������Qb�o��掦�cr8��|��Gx	٫j�2������V�Q8��rU��w�W�(-�/���E���=�@0��^AE�@��(�e�0����¨	0;�7o��0<\�� U0��\��5�!(���N���-�����PT�E�=�B|�*�Y��Y_�������h_�J�Gf2m���u�x'8 �l&.�
�V.�ɧ���\�)^ (-�ּ�������F���^Ed����O}��V3*:����w�"��l������\uW]U �	/,1� �S�Q]��b	x��M���R>h���9�KvWk��U@c����ۄ�y���Mqɓ���ˈ~L^TT4ΑO��[���-�ar���PQ�	@dlT�@�KE���fm�3|	i������x���T���;)�V�@�WP �a�H��!j�P����"���e9�Y��ɿ�e��JONK�G��j�Q��3[Ξ����z���� ��/Bh�&�"'�*6�e_[Ȣޅbƀf�r��O4{ ����ٖ�j�s�Wj�mZ`$a�G������$��p��#ڮ5��oϤ���$���&�s1m
�q�]�O�.��� ��ٳʿ��\��g�� ǯ���^���\�9P��X4�,�$��[N��E3 ���V��!\�Ҷ��*&uˢ�?w�4�A��,ּ����ݖO}�1ߑ��+,؀�|��͚����u��r`T����OV
.  ���Ѫ�u���\��o���|���^�#"U5ፗz8�H�(��g����,��^A,1jF���DZ<�<�0J�1	�7M\0���<V��ym{נ2ς�b��FF:sA��,)���,?��� �N��OӶB';�T[C�y,0�}[�&'���<��d�XHY��,��ZB�*(���+�7b6� u[��%r�6����~+wQ�d��f�ӷ��ʃ8,� �j�;78O'fK��, X�L�����C���?�E�nw~�"��#B}&�&?�0]C��d���']�q�1����V �^{Zw��Ql����z�w��B:��(
,������!����'�Bl�
��e1�<���,�£���ַp �``�^�푆%�=,t-��nf~��R���"�K��9`�[��%4�v"����D�	i��ُ m�K�����N��~!PP52�F�v���r�5�FǢ���E�
O�H�pl b��F����5�@�f!x 	�Y ���fH����	��* G@S�b�-(v�ᒁ{R�?5%DDm؈����A���&3��[P��%@�Q�I�%�� �,�.Q(_��w *	c��EA)�k�>��S]��⊢?E���o=���2U�nOJ�+��z{H'=m
Lbʍ�E�؞�y���7S�P�A�n׉��k�\�-!���P%�D���S�� &�"&���_'}<��]1�$}�*�Aޖ�pi%�t$�$�b���>�,d�qEO$7H_U; '�ٽ�{]��5�7��+܀~�O½p�Y�W�p�/�#,m��Y++_�'4s�@����s��Cք��!F��KKS��޵F��S:�
������G�7��"�S���eEb��PD�Vpm�Ij��,�Zw�.��u?E�,�/E�d2g����L��-7�n���P�b'b�)�"pX��"�け�Ra[�̶�Gܼ��{۞� ��'��hP�ٓ|Gί��c�Sߦ�w!�n���5�/��f:�4�V/��#�٫!��]�?ձZ�['���� <��+�*K�K4��BJ�QQtfvfi��~Q�?���n�1�̜y��F�޸�&0~j���5%�.tp��`N:\Pvl��%��Np�U�r�".���%�R�1����Z�U,a��7m�_�����L��ۨ��̊>F��h�hK�OS@�UH�N��N�8��Gf5Qг�tY�&�I(ݳ��xm@����������Npf����t�6o(ż�PX̿)�Ǣ�|/A�@�����B��hy�'�7���_L���"�� ��D<�w���͎�>�`n�%�Z���p��}����uut,Ü<|�Ù�!zT6Z��Ӛ�XD��"F��Q�FA����B�=p�^��=�@�NN�ߗL����:��m��<��psԹ��;�v����0���;[�k��;��)of��H
oN���1@��3�<+����<�n�o �<��3�tͳ+n�����)����4������?h�ߔ�M��Ԕ���vi��49�����bn��N������:�<������m7%Ο������o��/M)�·��*50��p0�^c��^>
W}��{�C�����Х�.d�����"99٫jO)'xw{~����}������1��C?�#�,^~�<����	~�GUph��ck���ח.]o�̓�:5�}!��G��%���em�GS�SN���ܜ0V��Y��gZ(��gu$�T4�M��%>���]��9.��GA�}�h���v坾��YB{�v��W�B��c�������~cᨁrҡ�16�-���'�,��1��6MZ��{<������ڼ�Q�?���>ބ��?�3(�稷��N���x#������`�k�k�����8H���U393k��D�XL{���;t!�2��6��x�3��G�Y�͛����Д�n��w�4��O�%n3��J��|*�u��v�C��L�4y�}R�w�(�K���\��-�wԋ�&��tV6������Ŵ�OI2|1yO$A�|S}��7a1�x�W��,���Q�&�חx>#�
[�O�7a����.��df�I	�����͙S.ڟ��2��{2��X�ЩX?/���Us�J��bӝx"��?_�7����� O:�t�k�E�����|�}�R�D�~
�S���?
���(XL֋vށ]��~��%�����ze��N���3�C˿<DN�^~n�m"�u�o���2���ny������kGd��y��Ky7��?�J�����?���g��_<=�kk��ԄD8� �>�SQ�	?��E��uM#�\��}�� J������)����wZ�o��ۏK
��x����8r��Lv9#�+_��ZB�]��PP�m�ޡ���D�c`�������Ңh�)w�ܒZиvA�a�$�?�%���.d�W&����ʫj	�bX�y���ff�@�V#�$�X�eBƲ���Ft�T��1���NyJ�*%�N�>I����E0�^,&�}��?z�iwKEpt��� �q�l�3?<<�vtr*��= 0^�q	B��u����o�����.���r>����q7���,������7u,ڌO5������Q��c��/�P[�A���Q�d��HUB�?���t���*A������L]~;��wh�h���x\��ܼ}֔V�8��t'�Wj_XU�$!K�e����%/3V �˯;&��A�ǧ�6a1
y|�v���ڻy�~����n��sU�b��_�M/�iiq��"}��7˿ՠ]��[�8�ay�̕�Q�1�/�H�t>���!�Qj�Ӛ���}@���os�ip����2�Y��������F��>�n�Y(�Ï�Vp^���`@`FYoT"W-衆�`�����i{���x��r4-��9ދ]�rO�l�-���s&�����du]zެ?���z1���a꧂�"��I���~�d��2^RT]�n6s���zM-Ai]��#5|lGq�����r�^� N�(���#��ި�H0˝={���wI{Dy�d���Ӽ��#ɶ��%��^-a���l�J� ������8,�J�Em�6�n�DM�4�t̜�n��>�P��:�5m�����D�KА!�B����u�)�}-���T~=~��U�ߠ$���_L!��S�5i�%P0*t��G��D*e%:��E㪷���_�y�߾ ��BZS��&�/������tQh	�J^SVYЉ�k
���x5���ua������'�wp�1� �Ŵ�Gɤ�����.gXٗ��!:w�Y�[q�xϾ�W"���K�a`�u`��`�,�
%~��ؔ�6��_��+��_�~�~n���]�z�,//�9gi�hևf���,ֿ;.F�[sY��{z���B�I;SS�� {{�g��%�Ѵȥ눃�c^��q����o!^8...��˯�B�β�����;��F3_[��zG��Ƿ�]�G�ߓ#x����g�PЫ�0��#2zz���A�6�� �\���55���f.[�
zC���Z�#��`p'��9��a�1y���I��yMj�J�i_���N�[�p�g�g�-d�Z'jiWD��Y���Lr�r�z�Z}Uͧ�4��o���΋Q�/zc�'&&:B���a�����(-�}ݛi�ҕL���V8���3��i݂��v=ƀ��n7Xv$K��̉ϱ�U0V�ēL��V�EeƟ#�SA�Nv��֨&��5������N�|��/5�i�kwuԶ���ZV_��6Ô5x/|!b�;�F|�A��^Y���S4%��gS�A~0ӺX�4���=p�pi�=���0�����e&� �TO���t !�Y��t��i��$�LVv�qb��G��G�î�=�C� �>�lr��������|�4�F[�,���5w��yjTXT�vw�yvW�R�R��6����e�wvc@����NiM�`ɐ7q��IȆƞ��23�h���ր�f�����gr-�g�AU�9�aG�c ���+���v@��h1�ѝ��3��U=��H�S���!C�X*�9���/�Lc�@Y�&�X�W���U���I�}��ZZZB�
_s/vuV�f0P(�섩AV}z�y~y| Xk��7�͵Y�CXd�*䁣�YH���=}�`�55�J�@���ҫS�~S��I���U��č�y�<i��1�i^�;�g�5�5T�83.f��6М8����hݳݛ��5X)�<����L�t��q>}8,Z��5�kbi�^�CM@�ib��K�&�cl�܆��0d"M���f��ԅ�����V����V�2�u��+a鹝Ú�D��� �	����>9�o^���5X��������N�5���D��ּ;���6�*ÜU��0%��u��.�hfV^��?�)Us�ҥK�>-P����|+QQ*n��7c	�u4D���0��Q��Ty��h��Ma���j�_y���Ȟ�9�����?�%��X��%�ld
u��>����ߍ"�~�7�!Xs��8U�']�>�>��q3N�=3Ů�ג՚�'�P=wl�^�����xX߼�{T�߀.B}�$/slj�,�4y/=�L���E]K+`�L�e@NϚ��Ԯܤ�g�2G��t!�D>�^6p5^�_���~�2:�3Ͱur�]i�JN��N!�>�<�L���oAB�����&Cw��Q�2tْ�SX8������L���ʛ�6,�'6�]��q�t;�^7X%p��u6ͭ���HSd��/��b��q�:gz9Z,�[��l��w��MK�6�H-!�H��1:��؆��I+WK����)-���z)/l-T��f�l^�vIc���� �,�
�;у�� �&{�)N���5Qtu#�¢����X2�N}�gw!{H*++�}�}�A�@V�'C�<`<����3�JʾX�b����2=>��
_��d��B��>}���S��ѬQ��Ǥ!{�K���N��k��֣< �=��ƐH#G����).�ye�I�[����KQ�~�6q��S̵TI�M�	�����~	`� ��C��_Z��<{���Y �];�^mМ�(�JK}����`�X�E�p����m<w`h�U}�G�܁��Ԥ�;����-=== `�$��6��s�������s��}@�3=n�'�~���uX*`z�{
���2Q �^G����(���$,�F6B�#Ѐ����.C��5�EY��M����&|�U�I��)h𩏣pӄ�]��W�����Eݟ��W8����?�O��F4���A��(Ih������(7�.�2��P#���PY����2�׳�>l��W��!�F�ͽ�(��3�	��k��¦E]�_�~��u���+}��1\l�t^m��ҷ�(�䬲�1V�>�ϵ���n?{z��C��p�V�����7�Q�r+0��r��3����a&�9�rZ�OB;�c_c��H��-%y�w��߷�~Oc��AF
E�P�`=L�ꃶ��"�څ�N�0�Y��{���[��������m����n/ŷ:�ܱb����ML~%�pp������(��[�˺��Rʍ^8�Xi��Q�5��C��%�%^C�I�j(�@�J�12�������(�}���!��-k�K���mɟ��-��W�@�I�hF4hf���
�.�TT�C=��$��Q�ԀV�k��F�R� �}S�
� ���m1�f���V�t_�$
/A��Ð��9�L�)��n���[��IHJ~�G�]�g�ÈW��S�)���^{�OЃ���P����")3c�`A�tK[��T��/L�ϩ��p�rBMM-OE�P��1�҂�YF�6m�<3��z`}�rXߚe4�rQ�V}9��9�s
_uv/��j���Hp��ڂ����gA��c�jΙ"�2Q��UfM�����AG��e;x�(Q�~��*�6AD�Km"�']�̍���6fU��P݄�1�sz�d��k�5��@���j��=�U�dV�摻vU%@EWCĈLi��h�?�	7����2��
�V��1=�Ll�ѯ��V�ڲg��j��TR2�c�4Zw�<^�PqK�ak��O��>��ҟ�ּ�
����u�����e
2�'�l�$�4�?�9Y$ؔ ��VVF�8�Y��o�}�Xt��l2B��Tq|*�G�/Ͼ����K��5ss����.�ӌC�D���@��t�*[	��hǾ�|g��!�$�O^������I��W �,�$U�$��/����r��O�}��f�|v�g����Q�@�(�G��u�-Wj�������}��h�k�Ǧ\��{�� UN@�;�tkS����^U�L���O����
�f�ZWf^$�?
ι�b�
'N�;��'�Al���.�q:=F���߃fc9�KTϹ0\��t�ji���|�@�q�ӂ���;��s��� A��ck)��a~'Tɓ�پ�>}"_�@��bS&������1lT��W���XL�:�$���e�X��d�j)L�ٱ��}ך��2�!ٹ�1cu+��'i<����<�T��~�����i��lG� i�ް(���/���`���R&r��08g$*Ůt�L��w���� � ^�p�e��c,8?c�ax>�Pk�|%�*�&7��؜Q[��9�'�>���v�'�]��sI�Af�[���Db;��B>�px�I
I�k��q 7NE���%}�˯@�(\a�c+��Sؚ.R�A��}�"�/
��'���}�h!�Ѷs{�\ў�����2��ln�Z`=����h��
tғ6�Zq�$W�%��h���7����Ӛ/��)�%��צ����dZ�~{}c8�p`�K�]l�L�+�����"��~=��u� ��i��t���â�r�p�l�j��t��V$��R�~<�*�Ni�����® fMߋ�����׭���K��T+���O��Zd'c��-�	�����n��3��JNf}��kOk����m�n��-hj��hv�JY1iȍ���� ����S��5���{/�9�N�
�D-Qa��T<�\��ZF;&!!q<����-"��Ϛ�XL�cz:�A����B*Z�ZC[������{���l��#dZu8�0�D$�m=��e����k#�T��M"R�p�!R
p�z@<+>�xӍ��I⿽�h�H�H�f,ӹ^���S�h&@3�N� ��k��ӕ�'�[�9�	����@]���S�<p��x��^�1�/��/��K
�ӽ��'�)K	��7Z^�ӻ?�Oo��P\ʕ��n�̶�ї�Fo���+��O�Q�,sb��<]d}4c���A�p"ǄO�p3Lw�k]��LO�Y ���ȩnu
Db�S�!�~$�;NUM������n�Ѥ��/�b3@�<~���mڨ�6_E v�H���N�2�^�k�؇�?� r�6�F_g��ޝ|d!�:�5��bGbG�?lA4F���1�����u��4o8-��
���L���	��EsI�c�t����`�=z�ś������ϻA&���L���-���l�!���Lgf�^��ͼG=�e���I9U2��M����:�,(�|Q���.�[�a�ID�'͎��r�$�W�/]���]��j��fS�u�E���P%Mz�9�������l�N�.�Y8�q�\��U5�����0�s��&��_�?�N��^��&� 0��IS�|�6�7{��]��Z�d�N��k?55UJLz�j�Q�3~���1,#���E|�i!�H۠³y�ORAȞ�V̳�߃�LQ���U'ARކڦ�����p��kEH�@�m����+�zj���ܾ7�(�G�+8�C����ҪFE��>ݛt1ݣ*��� �Q��'��i���deHr��@V-�ܱ��z�Z��2�ո����Ya��E����Wt�P2�Rj����.��|���h��eT��r�&c����X����i.""�%^��ޝ�ƛ�H�A{~�6�3�g
�z����A�G�m�9<'����h�����-��YK,p��P7!��� S��{� >$�[�=c�㉤�bQ�o���+�x��TV�`��d�����	��(�u���vq&���2�+��Ϻ�h&⪨�ʞ������
�tO7j�xq��>�쏄8����u�k���~nE̋�y������ q�������J�DYFW��f7���~��s躛ڳ/��S7�J ��F�z,�B��Y�R����B��"?��\�j#���{=h�ǻ�i���d�Z�Md��IY���f��=�e[eJ���O$�h�Z�����3������g��?�=��d򀊺�ff���K<f�*p�юաVέc�ЃZ��|�;��a����4���ܢ���20�̜�~vY������N���!7�<�Q7�8��};"qޞ��>>����t3pX�8�R{��4OQj7L��xT3z�_�8�g���s u�h;Cy
�[�m7^�{cl|��#����}x��S��VE��.��<���B.�}��Jl֩Hs�\��Ɋ *Ԩh��BeB\�,UaD0���-��DkY�B�����s�{��T`i�v�?n�D>"z�	�8A&}\
��Rl�1�B�.H��� ǘ�6n3zp�/u�E�X
�bE�4��>��~�J�
cX�1�䞟���b��:�',@��s�z��1}WMЭе�9*>�)�=7�	t�3Ʌx	0���K�c�*Z;�#���}�
؎}�2�VW&Ϙ.ӭ8۷!��]��Q9�B�T*+N	����qjp���83W��ّ ~ϓC�/�Kr.�7��!�O�w�R�d�dq����}����&ɥrxɲ�h�УQܕVH}E���T�eLגIj2�zP��������v��l���
CI��"|,L�M����Lf�%p���6�Dg �w��5��0kɟ� �.C��@� A��
��)qk֥��"�$����jg�@��#y��I:4���Y�Ā� *2�ھ�^��� _\H��� ���j��U5���
#�61����� ��M&iI�2$�w`���V�I-�J�� �LR�����%$�Q�I��޵�`����<���NB���ND�0Z���ǭ�	d��n@�֏��I�k�͞�t�kW�g���Xu��_����j0�b��:�F�����K�4�#���T���mܯ�<x����#���2�`Ц����?Ae]@�����\�}�o�S���!G����
� r�����]܂Ԩ;T	,��6m�B^spO	ZY�m�n�, }�f�}	�{�H�w����ߖ������!����D��f/i�Z��b���f��(��ϗG�H����VAB��ln���%�?���뵸����@�b���9ovJ�N��䑞n�	���Ϋ��T�$}���� �W���܋e٤!�XI�B�H���S��ЃM�q%9inE&_��\��uF|�^�?�����i�'_�nuvH�+Ю0��X�.TA�B'� Ө5��H�"�VTTd�^$x��vŰl�;#�S��I����Cq]��jB�U��k�q��f�! ��t��wO��T����a2��Sa�v�k95]�`&�5�Ї1<�p�⹫���+���]�&�G�����B����{x�k�L���c�-�.*����[�X�RzC�����V�Nh���yQVƁ a
��b��ќ�b(�IG�pX��;�b������e�q�"٥�1mRh�ź�����,���eJ��h���%
���}�,���vq.�����q��wR�B�J�h4�	�}Z�WO[��)�Ľ[�� r��T�`1�8
��[��P�!�ֳ:�N}q.��J�OԘ"���C�:��H&E�}dlL6�y�E���������/pj�L{��s]T�m@O��rE�+�e:�bf��!���<��4�8oSm_;m�2Л�Ye�'�L�-�}'`{c��S�wyYp#��*j�*&�j�/�!��9WLw�l�S�� �1,� ��
3��j�$�Ǿ�c�SQ��-@��i�n"��%�_j�(3�N����xiKX�J;���`L��!hOv2������m333
��Ѹ�� ��8o,��]�Ӎ��]0�ڿt+�]�&����|��zt+z�74����J���h�G��� }L=�I�I��޵&�l�9i+Y]1�^:d�RTxhX�� ��lgr�t�z�Q��� y�����T��c�Z`���d�"�b�C�E���u��
�'*���N�TD�Oa�Q��!�t��?�S?͢t���u��g�Z$�E��f�'�橡�G ��w�X*�,'_�����a��u�p���B�2����-�O$rI��s��(j��DL����J���9�CN�E=����)���{,�`���B��
���g=;���w���K_?A��3��t����d�弐L�~7[b����畗CH�N�¥J5�ȋ&U�&�\\�&L�Pe���҈$X����4����?D�vi��U�4���!�APA�%a��
���	�q��+�"� Р� � F�$�������eWM�TMM��?4���}��s�Kr�<��ƠM��'2���=W��!������ku�X;u9ߠ �o�5:i����Ѭܢ"�)cSj�9p\#�z��o9�e��,�ވ::4T�*�$�'�������_�LhV�+��97>42�f)	uq�����`������2hP
AE������ӵX�9�\�`�ms�O'�To����.��K`�.֭�ov�B�5z���:47�����m��|�CRe�"-�G�4=8%L|h� )*�D�ۡ�r�Rhe-�"��"݁�	�333�����_���^�Ű6+�F� X�"���O���D�Ͼ��~i09`M�c��c���n)���4p���6i�u���KR���T��y^3u�AcڍB܅��s������C��{?}RO��O�s�h���P�e�W�As;'�U��T�n��Ƴ��<H'�it�t�;���X�;��t����Gտ���S���-Po:�w��\����I�o@3�9�ϟ�=�j�-�8+�)ڦyS�]�-��|dg�
v~1��|i`F�mJ��Fe)g��}� �4�~���L�X��5��x��-����XJ`���d�jO���b���&-D3P��I"~L��g4�vd]��o�(��Y�� nL~��'H*�;�������|��ZO����SÐ��*�E��u ���~�߇�
� �J(f���޵1I#���i��4w	�[7�:�ʬ��r��Խf2�q�!z|p��+"�Aޡ��'��Z]]��5���I��^}ceip(�����6r$�W�Y��C���i98=����i��~��Pcj���	��"�����b]��&�q+��b�G�;I�`�H��9֎�*��Z�E�����!�<�B]_�W��S�066vy~��i�_�6V�?�fИ�Zo��gǳa����(~� �RHP�����t*�\��$�t5��ѸKpX0�)�?��]֜[	�3L����7��|9�µ���_052�5���B&h�'�M��}η�N�b�Wśf�1j�f �C���Q),�DK��@	��g���^���M���*Ć;)p���v�u���P�,�\�s��^@��|�������k����###��'4F���G����~�Ih���b�ξ��2���n86��k]�(����=�N��m�7XgD�2{�^�*��-��<�}�W?��UaO�}���4T����ƿ�`X� ���l����KGڵ���&>��X�`;;a��\qE]�_oc/�A*�ŀ[	G����9(]#��w�V2p'�qP�;�h_�]�n�>\)<\W1[%�yҮ�hX���^#��Δ���A�{�;��p�v�-���֚h:��.����!�;0�*뤣����S�r������j&���V�w�^�	܊�U���\��@�o����܄,� �9�/5U��uu��v&��ָY\�t����W�#�l�a��gw��ЖR޳� ��+���l�h,|�7<	�Z�x�~~��O���G �k�~ɣ��AX/FjdEc�;�[>K������[���4+HC@�P)��Z���!��Y���*;�	�tPRw���[�|�����m��v�1>�F"5��0C�_g��2S���-��rK�☽ٔ�rIP��ל���9M�R p�@�n�ؿW�f��{�bF���Z���~:8���xI^����[�M w����!�W'�!���O琤��Ҽ-�s�3��S��|�.���
��g�NR�|;8�� ZOD��.��[�Ei��P:�k��=&,EͿ����5��(T����`����T�POiI�ͥ:��L#���� D`�V�&�+qde��U�1t52*w���� �E/�(�DO>�m�U� ��nS�°���R�6I�nC(��w��e��ޭ��3K�`�b���������}�0l��_��������t�jw�?�!���}C~���t�Ƙb��K���4�Ǻ���/:�3���vCq��'�.��7��p���m��+W59-�>0��æ�ˉ�r^�ƫ��䃶����I�P�����0�Έg���������f��?��{��j:z�o�[�.�V�#���aNat�4V����J��4�n��c�rg�Vl�� ?%�[�=(^�IƜ4� Wq������I,����[ 
���y� a�I��	���b�z׭f���+�CK�C���y���X��@�DvV���d�q�~{�4B#]"yټ�d���6�5\~3^�Ix�Y"2��i�0��GK6S�l�n4��:�E��L@P��d֬_�҃A3>j(�����1�}��İ�� �, �Z�~X��w'���hc4���(�{���_�U����\3���n�+aN�p�.��f��N�L���!g���.��3�\�5U��A�����deА��T.��~���D���͌���^,�����XY��f�����%�/R (*j��FW�Fs���`�=������l����3(#%`(tC�G)��\��lx"v?N_�V�9GP�X){rk�dq^fT��d���X>�c ��'X�0�Þ����fH5��e�3�H_��cT���R��ߓÌx�:��8����V#�����Eu��~��,��`��@0���n��[�^���m&�*l��~y֪�pp�������L<~��_�P?
xw��*�@nb�� 5-+��	x�\wO�+��g,�Rb���	
**���C�~���(�2����5��"c;��*����	C�#������`��P�	)_�Ic-��b�?���ک�j�ik� ;k�6�@kn4����Ϗa�,1�cb�1,���c��MZs�ʧU�ޜP4!^���w�Lԥ���q�}�ꕒ�/�[��0gDA!�p"{E�?��N�s2)�Q#��ɾ�}[��s[��ꩆ��id2�5QZ��,�,�����N�Th	�p����T�$`�Z��fs�e�P.�4�ɫ~���@/��nU����ۉL�E�se�F���7I��`,_���z��Uׂ�Rv�ZYQs���=�K�˄V�~�L�;��̊�����'CmY�"_C��w̆˷��	'�Qo���F���_����+,*��Q5�X5���Fw8�J�''&�� .켷�(�Q�	�,����9Ws;.W���1��K�9&5E�,�ј��}��{�wY���&~+���G�H!͹��>ju��+n�a4_�̄w�����s&�&��'��u�x�~���-���@0�[����Ɗ�5P:bJ�LfJD���d�n���T���N\r6�?z5fԾ����רg����W�P�0�/Ϙ"�u����x��v�M��Z$H���lBxtw�J�r���K�M��1��<�1�U855�B5�Ue�Q'�7��{c�~@�6��@f_M��;��nM�&i�[)JW~�2(��z�oO�����rB������ܢ�mB<�hѷs�o�?D�!�����DϪ3��Y
{Ҝ���������	��_C��۵(�[��$0�?	^��R�T�uj��>�M�?Do֭�oÍW���%;�?B�wxdY�lo�|qT3���5��]<�R�~��sq��,
��o]]��5H�W�'=��3�3�ڄ4h��.����TtQsmaw�N�/[�s�+�L콣���� E��R&g���I�?�NI�_m��OK�:Ύ����D�+�$�lHY�<<�菮�e '^�NO1��/V�0O"����yၫ {��٤R�د����<�K���~�t�A�W-�i�i�-e�F�t��ϑa+�Y��X�	H8ƟW���݇�B��ZG +�Y�8� 8ߪE�{�xn]�[+�����c!����ƙj+Ʊ½v��0F2j��9��q�y�F���ɣ8F��#&�[�)l)��\F'`�j�-==}�+���yCaa!g�]�l�3�\~�����#V��W��EEE���.�m�x�R���&�U���;�/�p(%7�%���ӺaY��RGH��K��m��K�4�芨M����O#�uz1�c��;3Ir�n�R�L5��rnr6,zwZ�����ɧ�s���ׄ��F,���mhh�aMԝ�-���fo4˲��U�{K�+,���[�B�fgg3�j�Ǚ��m�/��	�\�<<b;v��N�g��'�+%��"q+:�ӹ���L�Է���s�g;!j�]�s�C��������58Ty��}�_�j�Фo.��w�k%w�41�iM�V�n����զe]Fg��������#=!��"�]ᠡ��X�Z��/�.ۮ���m$��c������(Z
5_�Z��wu�}��ZQ�C��{�N�����r2�����P��fF~p(AES�'Jς`^���i!ƃ��?�%$r���+�R�� $%�����h��5���Ԭ+���P�w��=���C��t.���ּ�&6N�vUD�c>J0wʂ�M�Wg6}j,�f�|6�u
�͞:���"Ӱ�<�-�Nɯ;��N�%P<P��.�B��Z�-��Ѭ D�o����	��y��6��4�D��a�iC	�Ncp۝����J��8Дc��6���eV0D��؃�y�s�?�{����V|�h3�-���t�v���$��Ӝ���6��ey�����%���^�v�q��V��S޼y�֢ڰ��3o�i 
�@M��|�-�P���t*�����)����a\(:����NBb�H�)��w"DQ���s��jP��rwK��������%>�r��L��z0�F��6�y�|�Gz#�%hf�0�Y�FJ9�y��Ǖ�����z�ޮ�%<z�8��4��)��:�����-�Se(�w��r�ՓO]�D%�,�����mp�p�U{#�EE��Y'�}����3X�x�C-?�4M�s���᎗q�X�?*ydEZ�f���_, $��������E�*;׳�7��7�y���~~_�F����Sc����T�N ��� ����Ӿ>`�X���'������J��TU����&�������k���(����}�&9{�.�'PK   �	DX��x��  $     jsons/user_defined.json�Y�n�H�A� ��Z���or��16c������M��D*���A�3�M[��Ȧ(���l�OW7�T�*��ax2\/C�Ň4˃���C�̊�1Y�������O7�v^͝�~������^tv��^����pE�*��,�ûQ��t��Ijg�0fp9��'�c��)���&H'F�P��;�a��l���2�9sp�r�51����WH� ��T8�Ƌ��ߒ
�n�pb��'뼀�,?��bx�c����l�����lY�j�^y�,�q���9�u�}[�E���Z�,�Y�P,���߲�&����A����kQ�ɪ\���l��n�o�>N�?G�	��a�G��{vq��_QXڄ�`/�2����	+{��1����&��*☢��{a��<��d��iP� ���-��@u����(�ibF��I��ߤ���m�����	��6)E�����A����\"�M>�G����)���(�v:�öp��t@Ҥ��p��J��"��t8W�[������$-�6NZڒ�d_�x|�-IK��5qԖ��{��8j�cu��M�Q�U�Q���A�x��-y��D�Dڒ�xO�8�hK�=Q��b-�K�D����$/��uW���Mm� ��,����$�\3��q�S�0��vORj��[��(�E(Wٶt��ˍ���75�|�We�����Ĳr8��j+���b�x���%n�e����X��k{k]OlE��S�V�
�WKo
�wX����"�����"p�s{>P'm��\ξ8뾆�s�-�>}��E��D��s�ʺX��Ugqe��1�J"h�RBQ�0A�M�+Z��^�V�X�d�d�j�eT ���"!L>}�����P�Y�:��1l�����c#4c#�(k�g�+�۫��*^�+Ji����ƅ@3W��]��JK�?�f�R����(����x@)f�zW#-����i<ҷHIr�
�բ*�1+t׶��1Kt�Hm-�c�uG���.9fq�R�#==��ǖ��A�Z���r��S)�0�oަ�:[�r�����"<^��3�]B��"�F�s�8u�'$��m�~�rY�l�8�\� &+�aU���Z9���&�B!�&	�)��b\�_zw��P5�$�v��lQ1�YbE�4�=�
�7ݦU�����_�ưS#Fj��4�[���}G����c�%PЩ�$]tzȀ4�VY���1�w��|zc=���!a�eXf˕�]xM]�)i��*�zF����W��«.%A�@�aRp"��z����$���������P�a��.sn�0�'��=�ť�H��

q�2R ����$Mcv�a���z��Z�S�9�JVk��i�Zϰ����y�
DB�X@ J�M`R�P�A�r'O���iR�y��)�[��6<�r��:��ƌ	���� �R�痚C8�z�D�t�t��ׄ~]�aq�8��\�9L�UF\�|�����S�2o�B�SIPpV#I�B��fB�P�a�i�0e�� �e�����ْ�Z���Ͳ??;�(�L%UO���x�SUv}MG`��w��:���њ���ͧx��B�����}}��\�E��2qYEKU��-��������c��d�{(�:�6���]�yN:�)!��b9C�C��
K9WN;a���Jf�3I�Hĭf(�L g(fF�:P���ma�U(��i�����E�n��H�D����רhy���`K�Zk���)�-�!��Q^�P�$��99/�����*�XW�;5D�g���w|sno}����K����?�HU��{Ŵ�8�.f���jC��[a�Ǵ�c������i�gs����9_�Pk������&�� >#y��̙`|@8T�w�іCeØ XQn�>Z����?PK
   �	DX�v{,�'  L�                  cirkitFile.jsonPK
   �	DXG�~��  � /             �'  images/0739a1b1-a163-452a-a325-ab452d55b136.pngPK
   �	DXd��  �   /             ��  images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   �	DX�Ƚ׌  �  /             � images/9185dcb2-65ea-4de0-8d42-42cedb1b5634.pngPK
   �DX*�e#o� Į /             � images/957f05b2-baab-48fc-bd29-824c654b1c09.pngPK
   �	DX	��#u } /             t� images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   �DX��dI� �� /             �' images/aa7df784-6767-4817-a6e6-80fad30d0eaa.pngPK
   �	DX���7z  �  /             z� images/be8de2bb-09ef-440a-a2d8-19619bf9d0dd.pngPK
   �	DX$7h�!  �!  /             A� images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   �	DX$[��>  dy  /             �� images/d3938c88-0382-4189-a86f-3cd234ee676b.pngPK
   �	DXP��/�  ǽ  /             �7 images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   �	DX/0�m  `  /             � images/f42dd85b-579e-4617-aa27-44ea24c5d2de.pngPK
   �	DXF���?� Q� /             e images/f590943e-678c-44eb-a174-3243ba5f3820.pngPK
   �	DX��x��  $               �
 jsons/user_defined.jsonPK      �  ��
   